
module wb_slave ( CLK_I, RST_I, NRESET, .ADR_I({ADR_I_4, ADR_I_3, ADR_I_2}), 
    .DAT_I({DAT_I_31, DAT_I_30, DAT_I_29, DAT_I_28, DAT_I_27, DAT_I_26, 
        DAT_I_25, DAT_I_24, DAT_I_23, DAT_I_22, DAT_I_21, DAT_I_20, DAT_I_19, 
        DAT_I_18, DAT_I_17, DAT_I_16, DAT_I_15, DAT_I_14, DAT_I_13, DAT_I_12, 
        DAT_I_11, DAT_I_10, DAT_I_9, DAT_I_8, DAT_I_7, DAT_I_6, DAT_I_5, 
        DAT_I_4, DAT_I_3, DAT_I_2, DAT_I_1, DAT_I_0}), .DAT_O({DAT_O_31, 
        DAT_O_30, DAT_O_29, DAT_O_28, DAT_O_27, DAT_O_26, DAT_O_25, DAT_O_24, 
        DAT_O_23, DAT_O_22, DAT_O_21, DAT_O_20, DAT_O_19, DAT_O_18, DAT_O_17, 
        DAT_O_16, DAT_O_15, DAT_O_14, DAT_O_13, DAT_O_12, DAT_O_11, DAT_O_10, 
        DAT_O_9, DAT_O_8, DAT_O_7, DAT_O_6, DAT_O_5, DAT_O_4, DAT_O_3, DAT_O_2, 
        DAT_O_1, DAT_O_0}), .SEL_I({SEL_I_3, SEL_I_2, SEL_I_1, SEL_I_0}), WE_I, 
        STB_I, CYC_I, ACK_O, ERR_O, INTA_O, BL, CSL, VSL, HSL, PC, .CD({CD_1, 
        CD_0}), .VBL({VBL_1, VBL_0}), CBSW, VBSW, Ven, AVMP, ACMP, bsint_in, 
        hint_in, vint_in, luint_in, sint_in, .Thsync({Thsync_7, Thsync_6, 
        Thsync_5, Thsync_4, Thsync_3, Thsync_2, Thsync_1, Thsync_0}), 
    .Thgdel({Thgdel_7, Thgdel_6, Thgdel_5, Thgdel_4, Thgdel_3, Thgdel_2, 
        Thgdel_1, Thgdel_0}), .Thgate({Thgate_15, Thgate_14, Thgate_13, 
        Thgate_12, Thgate_11, Thgate_10, Thgate_9, Thgate_8, Thgate_7, 
        Thgate_6, Thgate_5, Thgate_4, Thgate_3, Thgate_2, Thgate_1, Thgate_0}), 
    .Thlen({Thlen_15, Thlen_14, Thlen_13, Thlen_12, Thlen_11, Thlen_10, 
        Thlen_9, Thlen_8, Thlen_7, Thlen_6, Thlen_5, Thlen_4, Thlen_3, Thlen_2, 
        Thlen_1, Thlen_0}), .Tvsync({Tvsync_7, Tvsync_6, Tvsync_5, Tvsync_4, 
        Tvsync_3, Tvsync_2, Tvsync_1, Tvsync_0}), .Tvgdel({Tvgdel_7, Tvgdel_6, 
        Tvgdel_5, Tvgdel_4, Tvgdel_3, Tvgdel_2, Tvgdel_1, Tvgdel_0}), 
    .Tvgate({Tvgate_15, Tvgate_14, Tvgate_13, Tvgate_12, Tvgate_11, Tvgate_10, 
        Tvgate_9, Tvgate_8, Tvgate_7, Tvgate_6, Tvgate_5, Tvgate_4, Tvgate_3, 
        Tvgate_2, Tvgate_1, Tvgate_0}), .Tvlen({Tvlen_15, Tvlen_14, Tvlen_13, 
        Tvlen_12, Tvlen_11, Tvlen_10, Tvlen_9, Tvlen_8, Tvlen_7, Tvlen_6, 
        Tvlen_5, Tvlen_4, Tvlen_3, Tvlen_2, Tvlen_1, Tvlen_0}), .VBARa({
        VBARa_31, VBARa_30, VBARa_29, VBARa_28, VBARa_27, VBARa_26, VBARa_25, 
        VBARa_24, VBARa_23, VBARa_22, VBARa_21, VBARa_20, VBARa_19, VBARa_18, 
        VBARa_17, VBARa_16, VBARa_15, VBARa_14, VBARa_13, VBARa_12, VBARa_11, 
        VBARa_10, VBARa_9, VBARa_8, VBARa_7, VBARa_6, VBARa_5, VBARa_4, 
        VBARa_3, VBARa_2}), .VBARb({VBARb_31, VBARb_30, VBARb_29, VBARb_28, 
        VBARb_27, VBARb_26, VBARb_25, VBARb_24, VBARb_23, VBARb_22, VBARb_21, 
        VBARb_20, VBARb_19, VBARb_18, VBARb_17, VBARb_16, VBARb_15, VBARb_14, 
        VBARb_13, VBARb_12, VBARb_11, VBARb_10, VBARb_9, VBARb_8, VBARb_7, 
        VBARb_6, VBARb_5, VBARb_4, VBARb_3, VBARb_2}), .CBAR({CBAR_31, CBAR_30, 
        CBAR_29, CBAR_28, CBAR_27, CBAR_26, CBAR_25, CBAR_24, CBAR_23, CBAR_22, 
        CBAR_21, CBAR_20, CBAR_19, CBAR_18, CBAR_17, CBAR_16, CBAR_15, CBAR_14, 
        CBAR_13, CBAR_12, CBAR_11}) );
  input CLK_I, RST_I, NRESET, ADR_I_4, ADR_I_3, ADR_I_2, DAT_I_31, DAT_I_30,
         DAT_I_29, DAT_I_28, DAT_I_27, DAT_I_26, DAT_I_25, DAT_I_24, DAT_I_23,
         DAT_I_22, DAT_I_21, DAT_I_20, DAT_I_19, DAT_I_18, DAT_I_17, DAT_I_16,
         DAT_I_15, DAT_I_14, DAT_I_13, DAT_I_12, DAT_I_11, DAT_I_10, DAT_I_9,
         DAT_I_8, DAT_I_7, DAT_I_6, DAT_I_5, DAT_I_4, DAT_I_3, DAT_I_2,
         DAT_I_1, DAT_I_0, SEL_I_3, SEL_I_2, SEL_I_1, SEL_I_0, WE_I, STB_I,
         CYC_I, AVMP, ACMP, bsint_in, hint_in, vint_in, luint_in, sint_in;
  output DAT_O_31, DAT_O_30, DAT_O_29, DAT_O_28, DAT_O_27, DAT_O_26, DAT_O_25,
         DAT_O_24, DAT_O_23, DAT_O_22, DAT_O_21, DAT_O_20, DAT_O_19, DAT_O_18,
         DAT_O_17, DAT_O_16, DAT_O_15, DAT_O_14, DAT_O_13, DAT_O_12, DAT_O_11,
         DAT_O_10, DAT_O_9, DAT_O_8, DAT_O_7, DAT_O_6, DAT_O_5, DAT_O_4,
         DAT_O_3, DAT_O_2, DAT_O_1, DAT_O_0, ACK_O, ERR_O, INTA_O, BL, CSL,
         VSL, HSL, PC, CD_1, CD_0, VBL_1, VBL_0, CBSW, VBSW, Ven, Thsync_7,
         Thsync_6, Thsync_5, Thsync_4, Thsync_3, Thsync_2, Thsync_1, Thsync_0,
         Thgdel_7, Thgdel_6, Thgdel_5, Thgdel_4, Thgdel_3, Thgdel_2, Thgdel_1,
         Thgdel_0, Thgate_15, Thgate_14, Thgate_13, Thgate_12, Thgate_11,
         Thgate_10, Thgate_9, Thgate_8, Thgate_7, Thgate_6, Thgate_5, Thgate_4,
         Thgate_3, Thgate_2, Thgate_1, Thgate_0, Thlen_15, Thlen_14, Thlen_13,
         Thlen_12, Thlen_11, Thlen_10, Thlen_9, Thlen_8, Thlen_7, Thlen_6,
         Thlen_5, Thlen_4, Thlen_3, Thlen_2, Thlen_1, Thlen_0, Tvsync_7,
         Tvsync_6, Tvsync_5, Tvsync_4, Tvsync_3, Tvsync_2, Tvsync_1, Tvsync_0,
         Tvgdel_7, Tvgdel_6, Tvgdel_5, Tvgdel_4, Tvgdel_3, Tvgdel_2, Tvgdel_1,
         Tvgdel_0, Tvgate_15, Tvgate_14, Tvgate_13, Tvgate_12, Tvgate_11,
         Tvgate_10, Tvgate_9, Tvgate_8, Tvgate_7, Tvgate_6, Tvgate_5, Tvgate_4,
         Tvgate_3, Tvgate_2, Tvgate_1, Tvgate_0, Tvlen_15, Tvlen_14, Tvlen_13,
         Tvlen_12, Tvlen_11, Tvlen_10, Tvlen_9, Tvlen_8, Tvlen_7, Tvlen_6,
         Tvlen_5, Tvlen_4, Tvlen_3, Tvlen_2, Tvlen_1, Tvlen_0, VBARa_31,
         VBARa_30, VBARa_29, VBARa_28, VBARa_27, VBARa_26, VBARa_25, VBARa_24,
         VBARa_23, VBARa_22, VBARa_21, VBARa_20, VBARa_19, VBARa_18, VBARa_17,
         VBARa_16, VBARa_15, VBARa_14, VBARa_13, VBARa_12, VBARa_11, VBARa_10,
         VBARa_9, VBARa_8, VBARa_7, VBARa_6, VBARa_5, VBARa_4, VBARa_3,
         VBARa_2, VBARb_31, VBARb_30, VBARb_29, VBARb_28, VBARb_27, VBARb_26,
         VBARb_25, VBARb_24, VBARb_23, VBARb_22, VBARb_21, VBARb_20, VBARb_19,
         VBARb_18, VBARb_17, VBARb_16, VBARb_15, VBARb_14, VBARb_13, VBARb_12,
         VBARb_11, VBARb_10, VBARb_9, VBARb_8, VBARb_7, VBARb_6, VBARb_5,
         VBARb_4, VBARb_3, VBARb_2, CBAR_31, CBAR_30, CBAR_29, CBAR_28,
         CBAR_27, CBAR_26, CBAR_25, CBAR_24, CBAR_23, CBAR_22, CBAR_21,
         CBAR_20, CBAR_19, CBAR_18, CBAR_17, CBAR_16, CBAR_15, CBAR_14,
         CBAR_13, CBAR_12, CBAR_11;
  wire   ctrl_31, ctrl_30, ctrl_29, ctrl_28, ctrl_27, ctrl_26, ctrl_25,
         ctrl_24, ctrl_23, ctrl_22, ctrl_21, ctrl_20, ctrl_19, ctrl_18,
         ctrl_17, ctrl_16, ctrl_6_1, ctrl_3_1, ctrl_2_1, ctrl_1_1, stat_17,
         stat_16, stat_6, stat_5, stat_4, stat_1, stat_0, N66, N67, N68, N69,
         N70, n33, n34, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323;

  OAI212 U102 ( .A(n109), .B(n314), .C(stat_6), .Q(n112) );
  OAI212 U104 ( .A(n109), .B(n315), .C(stat_5), .Q(n113) );
  OAI212 U106 ( .A(n109), .B(n316), .C(stat_4), .Q(n114) );
  OAI212 U108 ( .A(n109), .B(n317), .C(stat_1), .Q(n115) );
  OAI212 U110 ( .A(n109), .B(n318), .C(stat_0), .Q(n116) );
  DFC3 stat_reg_17 ( .D(n268), .C(CLK_I), .RN(n62), .Q(stat_17) );
  DFC3 stat_reg_16 ( .D(n269), .C(CLK_I), .RN(n62), .Q(stat_16) );
  DFC3 stat_reg_6 ( .D(N70), .C(CLK_I), .RN(n62), .Q(stat_6) );
  DFC3 stat_reg_5 ( .D(N69), .C(CLK_I), .RN(n62), .Q(stat_5) );
  DFC3 stat_reg_4 ( .D(N68), .C(CLK_I), .RN(n62), .Q(stat_4) );
  DFC3 stat_reg_1 ( .D(N67), .C(CLK_I), .RN(n62), .Q(stat_1) );
  DFC3 stat_reg_0 ( .D(N66), .C(CLK_I), .RN(n62), .Q(stat_0) );
  DFEC1 ctrl_reg_27 ( .D(n298), .E(n8), .C(CLK_I), .RN(n257), .Q(ctrl_27) );
  DFEC1 ctrl_reg_26 ( .D(n297), .E(n8), .C(CLK_I), .RN(n257), .Q(ctrl_26) );
  DFEC1 ctrl_reg_25 ( .D(n296), .E(n8), .C(CLK_I), .RN(n257), .Q(ctrl_25) );
  DFEC1 ctrl_reg_24 ( .D(n295), .E(n8), .C(CLK_I), .RN(n257), .Q(ctrl_24) );
  DFEC1 ctrl_reg_23 ( .D(n294), .E(n8), .C(CLK_I), .RN(n257), .Q(ctrl_23) );
  DFEC1 ctrl_reg_22 ( .D(n293), .E(n8), .C(CLK_I), .RN(n257), .Q(ctrl_22) );
  DFEC1 ctrl_reg_21 ( .D(n292), .E(n8), .C(CLK_I), .RN(n257), .Q(ctrl_21) );
  DFEC1 ctrl_reg_20 ( .D(n291), .E(n7), .C(CLK_I), .RN(n257), .Q(ctrl_20) );
  DFEC1 ctrl_reg_19 ( .D(n290), .E(n7), .C(CLK_I), .RN(n258), .Q(ctrl_19) );
  DFEC1 ctrl_reg_18 ( .D(n289), .E(n7), .C(CLK_I), .RN(n258), .Q(ctrl_18) );
  DFEC1 ctrl_reg_6 ( .D(n277), .E(n5), .C(CLK_I), .RN(n259), .Q(ctrl_6_1) );
  DFEC1 VBARa_reg_9 ( .D(n280), .E(n26), .C(CLK_I), .RN(n250), .Q(VBARa_9) );
  DFEC1 VBARa_reg_8 ( .D(n279), .E(n25), .C(CLK_I), .RN(n251), .Q(VBARa_8) );
  DFEC1 VBARa_reg_7 ( .D(n278), .E(n25), .C(CLK_I), .RN(n251), .Q(VBARa_7) );
  DFEC1 VBARa_reg_6 ( .D(n277), .E(n25), .C(CLK_I), .RN(n251), .Q(VBARa_6) );
  DFEC1 VBARa_reg_5 ( .D(n276), .E(n25), .C(CLK_I), .RN(n251), .Q(VBARa_5) );
  DFEC1 VBARa_reg_4 ( .D(n275), .E(n25), .C(CLK_I), .RN(n251), .Q(VBARa_4) );
  DFEC1 VBARa_reg_3 ( .D(n274), .E(n25), .C(CLK_I), .RN(n251), .Q(VBARa_3) );
  DFEC1 VBARa_reg_2 ( .D(n273), .E(n25), .C(CLK_I), .RN(n251), .Q(VBARa_2) );
  DFEC1 VBARb_reg_29 ( .D(n300), .E(n35), .C(CLK_I), .RN(n251), .Q(VBARb_29)
         );
  DFEC1 VBARb_reg_28 ( .D(n299), .E(n35), .C(CLK_I), .RN(n252), .Q(VBARb_28)
         );
  DFEC1 VBARb_reg_27 ( .D(n298), .E(n35), .C(CLK_I), .RN(n252), .Q(VBARb_27)
         );
  DFEC1 VBARb_reg_26 ( .D(n297), .E(n35), .C(CLK_I), .RN(n252), .Q(VBARb_26)
         );
  DFEC1 VBARb_reg_25 ( .D(n296), .E(n35), .C(CLK_I), .RN(n252), .Q(VBARb_25)
         );
  DFEC1 VBARb_reg_24 ( .D(n295), .E(n35), .C(CLK_I), .RN(n252), .Q(VBARb_24)
         );
  DFEC1 VBARb_reg_23 ( .D(n294), .E(n35), .C(CLK_I), .RN(n252), .Q(VBARb_23)
         );
  DFEC1 VBARb_reg_22 ( .D(n293), .E(n32), .C(CLK_I), .RN(n252), .Q(VBARb_22)
         );
  DFEC1 VBARb_reg_21 ( .D(n292), .E(n32), .C(CLK_I), .RN(n252), .Q(VBARb_21)
         );
  DFEC1 VBARb_reg_20 ( .D(n291), .E(n32), .C(CLK_I), .RN(n252), .Q(VBARb_20)
         );
  DFEC1 VBARb_reg_19 ( .D(n290), .E(n32), .C(CLK_I), .RN(n252), .Q(VBARb_19)
         );
  DFEC1 VBARb_reg_18 ( .D(n289), .E(n32), .C(CLK_I), .RN(n253), .Q(VBARb_18)
         );
  DFEC1 VBARb_reg_17 ( .D(n288), .E(n32), .C(CLK_I), .RN(n253), .Q(VBARb_17)
         );
  DFEC1 VBARb_reg_16 ( .D(n287), .E(n32), .C(CLK_I), .RN(n253), .Q(VBARb_16)
         );
  DFEC1 VBARb_reg_15 ( .D(n286), .E(n31), .C(CLK_I), .RN(n253), .Q(VBARb_15)
         );
  DFEC1 VBARb_reg_14 ( .D(n285), .E(n31), .C(CLK_I), .RN(n253), .Q(VBARb_14)
         );
  DFEC1 VBARb_reg_13 ( .D(n284), .E(n31), .C(CLK_I), .RN(n253), .Q(VBARb_13)
         );
  DFEC1 VBARb_reg_12 ( .D(n283), .E(n31), .C(CLK_I), .RN(n253), .Q(VBARb_12)
         );
  DFEC1 VBARb_reg_11 ( .D(n282), .E(n31), .C(CLK_I), .RN(n253), .Q(VBARb_11)
         );
  DFEC1 VBARb_reg_10 ( .D(n281), .E(n31), .C(CLK_I), .RN(n253), .Q(VBARb_10)
         );
  DFEC1 ctrl_reg_9 ( .D(n280), .E(n6), .C(CLK_I), .RN(n259), .Q(CD_0) );
  DFEC1 ctrl_reg_8 ( .D(n279), .E(n6), .C(CLK_I), .RN(n259), .Q(VBL_1) );
  DFEC1 ctrl_reg_7 ( .D(n278), .E(n6), .C(CLK_I), .RN(n259), .Q(VBL_0) );
  DFEC1 ctrl_reg_5 ( .D(n276), .E(n5), .C(CLK_I), .RN(n259), .Q(CBSW) );
  DFEC1 ctrl_reg_4 ( .D(n275), .E(n5), .C(CLK_I), .RN(n259), .Q(VBSW) );
  DFEC1 ctrl_reg_17 ( .D(n288), .E(n7), .C(CLK_I), .RN(n258), .Q(ctrl_17) );
  DFEC1 ctrl_reg_16 ( .D(n287), .E(n7), .C(CLK_I), .RN(n258), .Q(ctrl_16) );
  DFEC1 htim_reg_1 ( .D(n272), .E(n10), .C(CLK_I), .RN(n254), .Q(Thgate_1), 
        .QN(n33) );
  DFEC1 htim_reg_0 ( .D(n271), .E(n10), .C(CLK_I), .RN(n254), .Q(Thgate_0), 
        .QN(n34) );
  DFEC1 VBARa_reg_13 ( .D(n284), .E(n26), .C(CLK_I), .RN(n250), .Q(VBARa_13)
         );
  DFEC1 VBARa_reg_12 ( .D(n283), .E(n26), .C(CLK_I), .RN(n250), .Q(VBARa_12)
         );
  DFEC1 VBARa_reg_11 ( .D(n282), .E(n26), .C(CLK_I), .RN(n250), .Q(VBARa_11)
         );
  DFEC1 VBARa_reg_10 ( .D(n281), .E(n26), .C(CLK_I), .RN(n250), .Q(VBARa_10)
         );
  DFEC1 VBARb_reg_9 ( .D(n280), .E(n31), .C(CLK_I), .RN(n253), .Q(VBARb_9) );
  DFEC1 VBARb_reg_8 ( .D(n279), .E(n30), .C(CLK_I), .RN(n254), .Q(VBARb_8) );
  DFEC1 VBARb_reg_7 ( .D(n278), .E(n30), .C(CLK_I), .RN(n254), .Q(VBARb_7) );
  DFEC1 VBARb_reg_6 ( .D(n277), .E(n30), .C(CLK_I), .RN(n254), .Q(VBARb_6) );
  DFEC1 VBARb_reg_5 ( .D(n276), .E(n30), .C(CLK_I), .RN(n254), .Q(VBARb_5) );
  DFEC1 VBARb_reg_4 ( .D(n275), .E(n30), .C(CLK_I), .RN(n254), .Q(VBARb_4) );
  DFEC1 VBARb_reg_3 ( .D(n274), .E(n30), .C(CLK_I), .RN(n254), .Q(VBARb_3) );
  DFEC1 VBARb_reg_2 ( .D(n273), .E(n30), .C(CLK_I), .RN(n254), .Q(VBARb_2) );
  DFEC1 ctrl_reg_11 ( .D(n282), .E(n6), .C(CLK_I), .RN(n258), .Q(PC) );
  DFEC1 ctrl_reg_10 ( .D(n281), .E(n6), .C(CLK_I), .RN(n258), .Q(CD_1) );
  DFEC1 ctrl_reg_2 ( .D(n273), .E(n5), .C(CLK_I), .RN(n259), .Q(ctrl_2_1) );
  DFEC1 vtim_reg_27 ( .D(n298), .E(n18), .C(CLK_I), .RN(n263), .Q(Tvsync_3) );
  DFEC1 vtim_reg_26 ( .D(n297), .E(n18), .C(CLK_I), .RN(n263), .Q(Tvsync_2) );
  DFEC1 vtim_reg_25 ( .D(n296), .E(n18), .C(CLK_I), .RN(n263), .Q(Tvsync_1) );
  DFEC1 vtim_reg_24 ( .D(n295), .E(n18), .C(CLK_I), .RN(n263), .Q(Tvsync_0) );
  DFEC1 vtim_reg_23 ( .D(n294), .E(n18), .C(CLK_I), .RN(n263), .Q(Tvgdel_7) );
  DFEC1 vtim_reg_22 ( .D(n293), .E(n18), .C(CLK_I), .RN(n264), .Q(Tvgdel_6) );
  DFEC1 vtim_reg_21 ( .D(n292), .E(n18), .C(CLK_I), .RN(n264), .Q(Tvgdel_5) );
  DFEC1 vtim_reg_20 ( .D(n291), .E(n17), .C(CLK_I), .RN(n264), .Q(Tvgdel_4) );
  DFEC1 vtim_reg_19 ( .D(n290), .E(n17), .C(CLK_I), .RN(n264), .Q(Tvgdel_3) );
  DFEC1 vtim_reg_18 ( .D(n289), .E(n17), .C(CLK_I), .RN(n264), .Q(Tvgdel_2) );
  DFEC1 vtim_reg_17 ( .D(n288), .E(n17), .C(CLK_I), .RN(n264), .Q(Tvgdel_1) );
  DFEC1 vtim_reg_16 ( .D(n287), .E(n17), .C(CLK_I), .RN(n264), .Q(Tvgdel_0) );
  DFEC1 hvlen_reg_9 ( .D(n280), .E(n21), .C(CLK_I), .RN(n247), .Q(Tvlen_9) );
  DFEC1 hvlen_reg_8 ( .D(n279), .E(n21), .C(CLK_I), .RN(n247), .Q(Tvlen_8) );
  DFEC1 hvlen_reg_7 ( .D(n278), .E(n21), .C(CLK_I), .RN(n247), .Q(Tvlen_7) );
  DFEC1 hvlen_reg_6 ( .D(n277), .E(n20), .C(CLK_I), .RN(n247), .Q(Tvlen_6) );
  DFEC1 hvlen_reg_5 ( .D(n276), .E(n20), .C(CLK_I), .RN(n248), .Q(Tvlen_5) );
  DFEC1 hvlen_reg_4 ( .D(n275), .E(n20), .C(CLK_I), .RN(n248), .Q(Tvlen_4) );
  DFEC1 hvlen_reg_3 ( .D(n274), .E(n20), .C(CLK_I), .RN(n248), .Q(Tvlen_3) );
  DFEC1 hvlen_reg_2 ( .D(n273), .E(n20), .C(CLK_I), .RN(n248), .Q(Tvlen_2) );
  DFEC1 hvlen_reg_1 ( .D(n272), .E(n20), .C(CLK_I), .RN(n248), .Q(Tvlen_1) );
  DFEC1 hvlen_reg_0 ( .D(n271), .E(n20), .C(CLK_I), .RN(n248), .Q(Tvlen_0) );
  DFEC1 htim_reg_27 ( .D(n298), .E(n13), .C(CLK_I), .RN(n260), .Q(Thsync_3) );
  DFEC1 htim_reg_26 ( .D(n297), .E(n13), .C(CLK_I), .RN(n260), .Q(Thsync_2) );
  DFEC1 htim_reg_25 ( .D(n296), .E(n13), .C(CLK_I), .RN(n260), .Q(Thsync_1) );
  DFEC1 htim_reg_24 ( .D(n295), .E(n13), .C(CLK_I), .RN(n260), .Q(Thsync_0) );
  DFEC1 htim_reg_23 ( .D(n294), .E(n13), .C(CLK_I), .RN(n260), .Q(Thgdel_7) );
  DFEC1 htim_reg_22 ( .D(n293), .E(n13), .C(CLK_I), .RN(n261), .Q(Thgdel_6) );
  DFEC1 htim_reg_21 ( .D(n292), .E(n13), .C(CLK_I), .RN(n261), .Q(Thgdel_5) );
  DFEC1 htim_reg_20 ( .D(n291), .E(n12), .C(CLK_I), .RN(n261), .Q(Thgdel_4) );
  DFEC1 htim_reg_19 ( .D(n290), .E(n12), .C(CLK_I), .RN(n261), .Q(Thgdel_3) );
  DFEC1 htim_reg_18 ( .D(n289), .E(n12), .C(CLK_I), .RN(n261), .Q(Thgdel_2) );
  DFEC1 htim_reg_17 ( .D(n288), .E(n12), .C(CLK_I), .RN(n261), .Q(Thgdel_1) );
  DFEC1 htim_reg_16 ( .D(n287), .E(n12), .C(CLK_I), .RN(n261), .Q(Thgdel_0) );
  DFEC1 hvlen_reg_27 ( .D(n298), .E(n23), .C(CLK_I), .RN(n245), .Q(Thlen_11)
         );
  DFEC1 hvlen_reg_26 ( .D(n297), .E(n23), .C(CLK_I), .RN(n245), .Q(Thlen_10)
         );
  DFEC1 hvlen_reg_25 ( .D(n296), .E(n23), .C(CLK_I), .RN(n246), .Q(Thlen_9) );
  DFEC1 hvlen_reg_24 ( .D(n295), .E(n23), .C(CLK_I), .RN(n246), .Q(Thlen_8) );
  DFEC1 hvlen_reg_23 ( .D(n294), .E(n23), .C(CLK_I), .RN(n246), .Q(Thlen_7) );
  DFEC1 hvlen_reg_22 ( .D(n293), .E(n23), .C(CLK_I), .RN(n246), .Q(Thlen_6) );
  DFEC1 hvlen_reg_21 ( .D(n292), .E(n23), .C(CLK_I), .RN(n246), .Q(Thlen_5) );
  DFEC1 hvlen_reg_20 ( .D(n291), .E(n22), .C(CLK_I), .RN(n246), .Q(Thlen_4) );
  DFEC1 hvlen_reg_19 ( .D(n290), .E(n22), .C(CLK_I), .RN(n246), .Q(Thlen_3) );
  DFEC1 hvlen_reg_18 ( .D(n289), .E(n22), .C(CLK_I), .RN(n246), .Q(Thlen_2) );
  DFEC1 hvlen_reg_17 ( .D(n288), .E(n22), .C(CLK_I), .RN(n246), .Q(Thlen_1) );
  DFEC1 hvlen_reg_16 ( .D(n287), .E(n22), .C(CLK_I), .RN(n246), .Q(Thlen_0) );
  DFEC1 hvlen_reg_15 ( .D(n286), .E(n22), .C(CLK_I), .RN(n247), .Q(Tvlen_15)
         );
  DFEC1 hvlen_reg_14 ( .D(n285), .E(n22), .C(CLK_I), .RN(n247), .Q(Tvlen_14)
         );
  DFEC1 hvlen_reg_13 ( .D(n284), .E(n21), .C(CLK_I), .RN(n247), .Q(Tvlen_13)
         );
  DFEC1 hvlen_reg_12 ( .D(n283), .E(n21), .C(CLK_I), .RN(n247), .Q(Tvlen_12)
         );
  DFEC1 hvlen_reg_11 ( .D(n282), .E(n21), .C(CLK_I), .RN(n247), .Q(Tvlen_11)
         );
  DFEC1 hvlen_reg_10 ( .D(n281), .E(n21), .C(CLK_I), .RN(n247), .Q(Tvlen_10)
         );
  DFEC1 ctrl_reg_3 ( .D(n274), .E(n5), .C(CLK_I), .RN(n259), .Q(ctrl_3_1) );
  DFEC1 ctrl_reg_1 ( .D(n272), .E(n5), .C(CLK_I), .RN(n259), .Q(ctrl_1_1) );
  DFEC1 ctrl_reg_0 ( .D(n271), .E(n5), .C(CLK_I), .RN(n259), .Q(Ven) );
  DFEC1 htim_reg_6 ( .D(n277), .E(n10), .C(CLK_I), .RN(n262), .Q(Thgate_6) );
  DFEC1 htim_reg_5 ( .D(n276), .E(n10), .C(CLK_I), .RN(n262), .Q(Thgate_5) );
  DFEC1 htim_reg_4 ( .D(n275), .E(n10), .C(CLK_I), .RN(n262), .Q(Thgate_4) );
  DFEC1 vtim_reg_15 ( .D(n286), .E(n17), .C(CLK_I), .RN(n264), .Q(Tvgate_15)
         );
  DFEC1 vtim_reg_14 ( .D(n285), .E(n17), .C(CLK_I), .RN(n264), .Q(Tvgate_14)
         );
  DFEC1 vtim_reg_13 ( .D(n284), .E(n16), .C(CLK_I), .RN(n264), .Q(Tvgate_13)
         );
  DFEC1 vtim_reg_12 ( .D(n283), .E(n16), .C(CLK_I), .RN(n59), .Q(Tvgate_12) );
  DFEC1 vtim_reg_11 ( .D(n282), .E(n16), .C(CLK_I), .RN(n61), .Q(Tvgate_11) );
  DFEC1 vtim_reg_10 ( .D(n281), .E(n16), .C(CLK_I), .RN(n60), .Q(Tvgate_10) );
  DFEC1 htim_reg_15 ( .D(n286), .E(n12), .C(CLK_I), .RN(n261), .Q(Thgate_15)
         );
  DFEC1 htim_reg_14 ( .D(n285), .E(n12), .C(CLK_I), .RN(n261), .Q(Thgate_14)
         );
  DFEC1 htim_reg_13 ( .D(n284), .E(n11), .C(CLK_I), .RN(n261), .Q(Thgate_13)
         );
  DFEC1 htim_reg_12 ( .D(n283), .E(n11), .C(CLK_I), .RN(n262), .Q(Thgate_12)
         );
  DFEC1 htim_reg_11 ( .D(n282), .E(n11), .C(CLK_I), .RN(n262), .Q(Thgate_11)
         );
  DFEC1 htim_reg_10 ( .D(n281), .E(n11), .C(CLK_I), .RN(n262), .Q(Thgate_10)
         );
  DFEC1 vtim_reg_9 ( .D(n280), .E(n16), .C(CLK_I), .RN(n59), .Q(Tvgate_9) );
  DFEC1 vtim_reg_8 ( .D(n279), .E(n16), .C(CLK_I), .RN(n61), .Q(Tvgate_8) );
  DFEC1 vtim_reg_7 ( .D(n278), .E(n16), .C(CLK_I), .RN(n60), .Q(Tvgate_7) );
  DFEC1 vtim_reg_6 ( .D(n277), .E(n15), .C(CLK_I), .RN(n249), .Q(Tvgate_6) );
  DFEC1 vtim_reg_5 ( .D(n276), .E(n15), .C(CLK_I), .RN(n62), .Q(Tvgate_5) );
  DFEC1 vtim_reg_4 ( .D(n275), .E(n15), .C(CLK_I), .RN(n62), .Q(Tvgate_4) );
  DFEC1 vtim_reg_3 ( .D(n274), .E(n15), .C(CLK_I), .RN(n245), .Q(Tvgate_3) );
  DFEC1 vtim_reg_2 ( .D(n273), .E(n15), .C(CLK_I), .RN(n245), .Q(Tvgate_2) );
  DFEC1 vtim_reg_1 ( .D(n272), .E(n15), .C(CLK_I), .RN(n245), .Q(Tvgate_1) );
  DFEC1 vtim_reg_0 ( .D(n271), .E(n15), .C(CLK_I), .RN(n245), .Q(Tvgate_0) );
  DFEC1 htim_reg_9 ( .D(n280), .E(n11), .C(CLK_I), .RN(n262), .Q(Thgate_9) );
  DFEC1 htim_reg_8 ( .D(n279), .E(n11), .C(CLK_I), .RN(n262), .Q(Thgate_8) );
  DFEC1 htim_reg_7 ( .D(n278), .E(n11), .C(CLK_I), .RN(n262), .Q(Thgate_7) );
  DFEC1 htim_reg_3 ( .D(n274), .E(n10), .C(CLK_I), .RN(n262), .Q(Thgate_3) );
  DFEC1 htim_reg_2 ( .D(n273), .E(n10), .C(CLK_I), .RN(n263), .Q(Thgate_2) );
  DFEC1 ctrl_reg_15 ( .D(n286), .E(n7), .C(CLK_I), .RN(n258), .Q(BL) );
  DFEC1 ctrl_reg_14 ( .D(n285), .E(n7), .C(CLK_I), .RN(n258), .Q(CSL) );
  DFEC1 ctrl_reg_13 ( .D(n284), .E(n6), .C(CLK_I), .RN(n258), .Q(VSL) );
  DFEC1 ctrl_reg_12 ( .D(n283), .E(n6), .C(CLK_I), .RN(n258), .Q(HSL) );
  DFEC1 CBAR_reg_31 ( .D(n302), .E(n304), .C(CLK_I), .RN(n62), .Q(CBAR_31) );
  DFEC1 CBAR_reg_30 ( .D(n301), .E(n304), .C(CLK_I), .RN(n260), .Q(CBAR_30) );
  DFEC1 CBAR_reg_29 ( .D(n300), .E(n304), .C(CLK_I), .RN(n254), .Q(CBAR_29) );
  DFEC1 CBAR_reg_28 ( .D(n299), .E(n304), .C(CLK_I), .RN(n255), .Q(CBAR_28) );
  DFEC1 CBAR_reg_27 ( .D(n298), .E(n304), .C(CLK_I), .RN(n255), .Q(CBAR_27) );
  DFEC1 CBAR_reg_26 ( .D(n297), .E(n304), .C(CLK_I), .RN(n255), .Q(CBAR_26) );
  DFEC1 CBAR_reg_25 ( .D(n296), .E(n304), .C(CLK_I), .RN(n255), .Q(CBAR_25) );
  DFEC1 CBAR_reg_24 ( .D(n295), .E(n304), .C(CLK_I), .RN(n255), .Q(CBAR_24) );
  DFEC1 CBAR_reg_23 ( .D(n294), .E(n304), .C(CLK_I), .RN(n255), .Q(CBAR_23) );
  DFEC1 CBAR_reg_22 ( .D(n293), .E(n304), .C(CLK_I), .RN(n255), .Q(CBAR_22) );
  DFEC1 CBAR_reg_21 ( .D(n292), .E(n304), .C(CLK_I), .RN(n255), .Q(CBAR_21) );
  DFEC1 CBAR_reg_20 ( .D(n291), .E(n304), .C(CLK_I), .RN(n255), .Q(CBAR_20) );
  DFEC1 CBAR_reg_19 ( .D(n290), .E(n304), .C(CLK_I), .RN(n255), .Q(CBAR_19) );
  DFEC1 CBAR_reg_18 ( .D(n289), .E(n304), .C(CLK_I), .RN(n256), .Q(CBAR_18) );
  DFEC1 CBAR_reg_17 ( .D(n288), .E(n304), .C(CLK_I), .RN(n256), .Q(CBAR_17) );
  DFEC1 CBAR_reg_16 ( .D(n287), .E(n304), .C(CLK_I), .RN(n256), .Q(CBAR_16) );
  DFEC1 CBAR_reg_15 ( .D(n286), .E(n304), .C(CLK_I), .RN(n256), .Q(CBAR_15) );
  DFEC1 CBAR_reg_14 ( .D(n285), .E(n304), .C(CLK_I), .RN(n256), .Q(CBAR_14) );
  DFEC1 CBAR_reg_13 ( .D(n284), .E(n304), .C(CLK_I), .RN(n256), .Q(CBAR_13) );
  DFEC1 CBAR_reg_12 ( .D(n283), .E(n304), .C(CLK_I), .RN(n256), .Q(CBAR_12) );
  DFEC1 CBAR_reg_11 ( .D(n282), .E(n304), .C(CLK_I), .RN(n256), .Q(CBAR_11) );
  DFEC1 VBARa_reg_31 ( .D(n302), .E(n29), .C(CLK_I), .RN(n248), .Q(VBARa_31)
         );
  DFEC1 VBARa_reg_30 ( .D(n301), .E(n29), .C(CLK_I), .RN(n248), .Q(VBARa_30)
         );
  DFEC1 VBARb_reg_31 ( .D(n302), .E(n36), .C(CLK_I), .RN(n251), .Q(VBARb_31)
         );
  DFEC1 VBARb_reg_30 ( .D(n301), .E(n36), .C(CLK_I), .RN(n251), .Q(VBARb_30)
         );
  DFEC1 vtim_reg_31 ( .D(n302), .E(n19), .C(CLK_I), .RN(n263), .Q(Tvsync_7) );
  DFEC1 vtim_reg_30 ( .D(n301), .E(n19), .C(CLK_I), .RN(n263), .Q(Tvsync_6) );
  DFEC1 vtim_reg_29 ( .D(n300), .E(n19), .C(CLK_I), .RN(n263), .Q(Tvsync_5) );
  DFEC1 vtim_reg_28 ( .D(n299), .E(n19), .C(CLK_I), .RN(n263), .Q(Tvsync_4) );
  DFEC1 ctrl_reg_31 ( .D(n302), .E(n9), .C(CLK_I), .RN(n256), .Q(ctrl_31) );
  DFEC1 ctrl_reg_30 ( .D(n301), .E(n9), .C(CLK_I), .RN(n256), .Q(ctrl_30) );
  DFEC1 ctrl_reg_29 ( .D(n300), .E(n9), .C(CLK_I), .RN(n257), .Q(ctrl_29) );
  DFEC1 ctrl_reg_28 ( .D(n299), .E(n9), .C(CLK_I), .RN(n257), .Q(ctrl_28) );
  DFEC1 hvlen_reg_31 ( .D(n302), .E(n24), .C(CLK_I), .RN(n245), .Q(Thlen_15)
         );
  DFEC1 hvlen_reg_30 ( .D(n301), .E(n24), .C(CLK_I), .RN(n245), .Q(Thlen_14)
         );
  DFEC1 hvlen_reg_29 ( .D(n300), .E(n24), .C(CLK_I), .RN(n245), .Q(Thlen_13)
         );
  DFEC1 hvlen_reg_28 ( .D(n299), .E(n24), .C(CLK_I), .RN(n245), .Q(Thlen_12)
         );
  DFEC1 htim_reg_31 ( .D(n302), .E(n14), .C(CLK_I), .RN(n260), .Q(Thsync_7) );
  DFEC1 htim_reg_30 ( .D(n301), .E(n14), .C(CLK_I), .RN(n260), .Q(Thsync_6) );
  DFEC1 htim_reg_29 ( .D(n300), .E(n14), .C(CLK_I), .RN(n260), .Q(Thsync_5) );
  DFEC1 htim_reg_28 ( .D(n299), .E(n14), .C(CLK_I), .RN(n260), .Q(Thsync_4) );
  DFEC1 VBARa_reg_29 ( .D(n300), .E(n28), .C(CLK_I), .RN(n248), .Q(VBARa_29)
         );
  DFEC1 VBARa_reg_28 ( .D(n299), .E(n28), .C(CLK_I), .RN(n248), .Q(VBARa_28)
         );
  DFEC1 VBARa_reg_27 ( .D(n298), .E(n28), .C(CLK_I), .RN(n249), .Q(VBARa_27)
         );
  DFEC1 VBARa_reg_26 ( .D(n297), .E(n28), .C(CLK_I), .RN(n249), .Q(VBARa_26)
         );
  DFEC1 VBARa_reg_25 ( .D(n296), .E(n28), .C(CLK_I), .RN(n249), .Q(VBARa_25)
         );
  DFEC1 VBARa_reg_24 ( .D(n295), .E(n28), .C(CLK_I), .RN(n249), .Q(VBARa_24)
         );
  DFEC1 VBARa_reg_23 ( .D(n294), .E(n28), .C(CLK_I), .RN(n249), .Q(VBARa_23)
         );
  DFEC1 VBARa_reg_22 ( .D(n293), .E(n27), .C(CLK_I), .RN(n249), .Q(VBARa_22)
         );
  DFEC1 VBARa_reg_21 ( .D(n292), .E(n27), .C(CLK_I), .RN(n249), .Q(VBARa_21)
         );
  DFEC1 VBARa_reg_20 ( .D(n291), .E(n27), .C(CLK_I), .RN(n249), .Q(VBARa_20)
         );
  DFEC1 VBARa_reg_19 ( .D(n290), .E(n27), .C(CLK_I), .RN(n249), .Q(VBARa_19)
         );
  DFEC1 VBARa_reg_18 ( .D(n289), .E(n27), .C(CLK_I), .RN(n250), .Q(VBARa_18)
         );
  DFEC1 VBARa_reg_17 ( .D(n288), .E(n27), .C(CLK_I), .RN(n250), .Q(VBARa_17)
         );
  DFEC1 VBARa_reg_16 ( .D(n287), .E(n27), .C(CLK_I), .RN(n250), .Q(VBARa_16)
         );
  DFEC1 VBARa_reg_15 ( .D(n286), .E(n26), .C(CLK_I), .RN(n250), .Q(VBARa_15)
         );
  DFEC1 VBARa_reg_14 ( .D(n285), .E(n26), .C(CLK_I), .RN(n250), .Q(VBARa_14)
         );
  INV3 U3 ( .A(n1), .Q(n2) );
  BUF2 U4 ( .A(n51), .Q(n62) );
  BUF2 U5 ( .A(n54), .Q(n253) );
  BUF2 U6 ( .A(n53), .Q(n252) );
  BUF2 U7 ( .A(n53), .Q(n251) );
  BUF2 U8 ( .A(n53), .Q(n250) );
  BUF2 U9 ( .A(n52), .Q(n248) );
  BUF2 U10 ( .A(n52), .Q(n247) );
  BUF2 U11 ( .A(n51), .Q(n246) );
  BUF2 U12 ( .A(n51), .Q(n245) );
  BUF2 U13 ( .A(n52), .Q(n249) );
  BUF2 U14 ( .A(n57), .Q(n264) );
  BUF2 U15 ( .A(n57), .Q(n263) );
  BUF2 U16 ( .A(n57), .Q(n262) );
  BUF2 U17 ( .A(n56), .Q(n261) );
  BUF2 U18 ( .A(n56), .Q(n259) );
  BUF2 U19 ( .A(n55), .Q(n258) );
  BUF2 U20 ( .A(n55), .Q(n257) );
  BUF2 U21 ( .A(n55), .Q(n256) );
  BUF2 U22 ( .A(n54), .Q(n255) );
  BUF2 U23 ( .A(n56), .Q(n260) );
  BUF2 U24 ( .A(n54), .Q(n254) );
  INV3 U25 ( .A(n109), .Q(n320) );
  NOR31 U26 ( .A(n322), .B(n119), .C(n321), .Q(ACK_O) );
  BUF2 U27 ( .A(n106), .Q(n38) );
  BUF2 U28 ( .A(n106), .Q(n37) );
  INV3 U29 ( .A(n42), .Q(n40) );
  INV3 U30 ( .A(n42), .Q(n41) );
  BUF2 U31 ( .A(n100), .Q(n45) );
  BUF2 U32 ( .A(n94), .Q(n49) );
  BUF2 U33 ( .A(n102), .Q(n43) );
  BUF2 U34 ( .A(n96), .Q(n47) );
  INV3 U35 ( .A(n108), .Q(n1) );
  NOR31 U36 ( .A(n311), .B(n312), .C(n313), .Q(n108) );
  BUF2 U37 ( .A(n106), .Q(n39) );
  BUF2 U38 ( .A(n100), .Q(n46) );
  BUF2 U39 ( .A(n102), .Q(n44) );
  BUF2 U40 ( .A(n94), .Q(n50) );
  BUF2 U41 ( .A(n96), .Q(n48) );
  BUF2 U42 ( .A(n310), .Q(n30) );
  BUF2 U43 ( .A(n310), .Q(n31) );
  BUF2 U44 ( .A(n310), .Q(n32) );
  BUF2 U45 ( .A(n310), .Q(n35) );
  BUF2 U46 ( .A(n309), .Q(n25) );
  BUF2 U47 ( .A(n309), .Q(n26) );
  BUF2 U48 ( .A(n309), .Q(n27) );
  BUF2 U49 ( .A(n309), .Q(n28) );
  BUF2 U50 ( .A(n308), .Q(n20) );
  BUF2 U51 ( .A(n308), .Q(n21) );
  BUF2 U52 ( .A(n308), .Q(n22) );
  BUF2 U53 ( .A(n308), .Q(n23) );
  BUF2 U54 ( .A(n307), .Q(n15) );
  BUF2 U55 ( .A(n307), .Q(n16) );
  BUF2 U56 ( .A(n307), .Q(n17) );
  BUF2 U57 ( .A(n307), .Q(n18) );
  BUF2 U58 ( .A(n306), .Q(n11) );
  BUF2 U59 ( .A(n306), .Q(n12) );
  BUF2 U60 ( .A(n306), .Q(n13) );
  BUF2 U61 ( .A(n305), .Q(n5) );
  BUF2 U62 ( .A(n305), .Q(n6) );
  BUF2 U63 ( .A(n305), .Q(n7) );
  BUF2 U64 ( .A(n305), .Q(n8) );
  BUF2 U65 ( .A(n306), .Q(n10) );
  BUF2 U66 ( .A(n308), .Q(n24) );
  BUF2 U67 ( .A(n307), .Q(n19) );
  BUF2 U68 ( .A(n306), .Q(n14) );
  BUF2 U69 ( .A(n305), .Q(n9) );
  BUF2 U70 ( .A(n310), .Q(n36) );
  BUF2 U71 ( .A(n309), .Q(n29) );
  NOR31 U72 ( .A(n321), .B(n319), .C(n322), .Q(ERR_O) );
  INV3 U73 ( .A(n119), .Q(n319) );
  BUF2 U74 ( .A(n303), .Q(n3) );
  BUF2 U75 ( .A(n303), .Q(n4) );
  BUF2 U76 ( .A(n60), .Q(n53) );
  BUF2 U77 ( .A(n61), .Q(n52) );
  BUF2 U78 ( .A(n58), .Q(n57) );
  BUF2 U79 ( .A(n59), .Q(n55) );
  BUF2 U80 ( .A(n59), .Q(n56) );
  BUF2 U81 ( .A(n61), .Q(n51) );
  BUF2 U82 ( .A(n60), .Q(n54) );
  NOR31 U83 ( .A(ADR_I_3), .B(ADR_I_4), .C(n313), .Q(n124) );
  NAND41 U84 ( .A(SEL_I_3), .B(SEL_I_2), .C(SEL_I_1), .D(SEL_I_0), .Q(n119) );
  NOR31 U85 ( .A(ADR_I_2), .B(ADR_I_3), .C(n311), .Q(n100) );
  NOR31 U86 ( .A(n312), .B(ADR_I_2), .C(n311), .Q(n94) );
  NOR31 U87 ( .A(n312), .B(ADR_I_4), .C(n313), .Q(n102) );
  NOR31 U88 ( .A(n311), .B(ADR_I_3), .C(n313), .Q(n96) );
  NOR31 U89 ( .A(ADR_I_3), .B(ADR_I_4), .C(ADR_I_2), .Q(n106) );
  NAND22 U90 ( .A(WE_I), .B(ACK_O), .Q(n109) );
  NAND41 U91 ( .A(n213), .B(n214), .C(n215), .D(n216), .Q(DAT_O_16) );
  AOI221 U92 ( .A(CBAR_16), .B(n2), .C(VBARb_16), .D(n49), .Q(n216) );
  AOI221 U93 ( .A(VBARa_16), .B(n47), .C(Thlen_0), .D(n45), .Q(n215) );
  AOI221 U94 ( .A(Tvgdel_0), .B(n44), .C(Thgdel_0), .D(n40), .Q(n214) );
  NAND41 U95 ( .A(n209), .B(n210), .C(n211), .D(n212), .Q(DAT_O_17) );
  AOI221 U96 ( .A(CBAR_17), .B(n2), .C(VBARb_17), .D(n49), .Q(n212) );
  AOI221 U97 ( .A(VBARa_17), .B(n47), .C(Thlen_1), .D(n45), .Q(n211) );
  AOI221 U98 ( .A(stat_17), .B(n124), .C(ctrl_17), .D(n39), .Q(n209) );
  NAND41 U99 ( .A(n141), .B(n142), .C(n143), .D(n144), .Q(DAT_O_4) );
  NAND22 U100 ( .A(VBSW), .B(n37), .Q(n142) );
  AOI221 U101 ( .A(Tvlen_4), .B(n46), .C(Tvgate_4), .D(n43), .Q(n143) );
  AOI221 U103 ( .A(VBARb_4), .B(n49), .C(VBARa_4), .D(n48), .Q(n144) );
  NAND41 U105 ( .A(n137), .B(n138), .C(n139), .D(n140), .Q(DAT_O_5) );
  NAND22 U107 ( .A(CBSW), .B(n37), .Q(n138) );
  AOI221 U109 ( .A(VBARb_5), .B(n50), .C(VBARa_5), .D(n48), .Q(n140) );
  AOI221 U111 ( .A(Tvlen_5), .B(n46), .C(Tvgate_5), .D(n43), .Q(n139) );
  NAND41 U112 ( .A(n133), .B(n134), .C(n135), .D(n136), .Q(DAT_O_6) );
  NAND22 U113 ( .A(ctrl_6_1), .B(n37), .Q(n134) );
  AOI221 U114 ( .A(VBARb_6), .B(n50), .C(VBARa_6), .D(n47), .Q(n136) );
  AOI221 U115 ( .A(Tvlen_6), .B(n46), .C(Tvgate_6), .D(n43), .Q(n135) );
  NAND41 U116 ( .A(n229), .B(n230), .C(n231), .D(n232), .Q(DAT_O_12) );
  NAND22 U117 ( .A(HSL), .B(n39), .Q(n229) );
  AOI221 U118 ( .A(CBAR_12), .B(n2), .C(VBARb_12), .D(n49), .Q(n232) );
  AOI221 U119 ( .A(VBARa_12), .B(n48), .C(Tvlen_12), .D(n45), .Q(n231) );
  NAND41 U120 ( .A(n225), .B(n226), .C(n227), .D(n228), .Q(DAT_O_13) );
  NAND22 U121 ( .A(VSL), .B(n39), .Q(n225) );
  AOI221 U122 ( .A(CBAR_13), .B(n2), .C(VBARb_13), .D(n49), .Q(n228) );
  AOI221 U123 ( .A(VBARa_13), .B(n48), .C(Tvlen_13), .D(n45), .Q(n227) );
  NAND41 U124 ( .A(n221), .B(n222), .C(n223), .D(n224), .Q(DAT_O_14) );
  NAND22 U125 ( .A(CSL), .B(n38), .Q(n221) );
  AOI221 U126 ( .A(CBAR_14), .B(n2), .C(VBARb_14), .D(n49), .Q(n224) );
  AOI221 U127 ( .A(VBARa_14), .B(n48), .C(Tvlen_14), .D(n45), .Q(n223) );
  NAND41 U128 ( .A(n217), .B(n218), .C(n219), .D(n220), .Q(DAT_O_15) );
  NAND22 U129 ( .A(BL), .B(n38), .Q(n217) );
  AOI221 U130 ( .A(CBAR_15), .B(n108), .C(VBARb_15), .D(n49), .Q(n220) );
  AOI221 U131 ( .A(VBARa_15), .B(n47), .C(Tvlen_15), .D(n45), .Q(n219) );
  NAND41 U132 ( .A(n237), .B(n238), .C(n239), .D(n240), .Q(DAT_O_10) );
  NAND22 U133 ( .A(CD_1), .B(n37), .Q(n237) );
  AOI221 U134 ( .A(ACMP), .B(n2), .C(VBARb_10), .D(n50), .Q(n240) );
  AOI221 U135 ( .A(VBARa_10), .B(n47), .C(Tvlen_10), .D(n45), .Q(n239) );
  NAND41 U136 ( .A(n233), .B(n234), .C(n235), .D(n236), .Q(DAT_O_11) );
  NAND22 U137 ( .A(PC), .B(n38), .Q(n233) );
  AOI221 U138 ( .A(CBAR_11), .B(n108), .C(VBARb_11), .D(n49), .Q(n236) );
  AOI221 U139 ( .A(VBARa_11), .B(n48), .C(Tvlen_11), .D(n45), .Q(n235) );
  NAND41 U140 ( .A(n205), .B(n206), .C(n207), .D(n208), .Q(DAT_O_18) );
  NAND22 U141 ( .A(ctrl_18), .B(n38), .Q(n205) );
  AOI221 U142 ( .A(CBAR_18), .B(n2), .C(VBARb_18), .D(n49), .Q(n208) );
  AOI221 U143 ( .A(VBARa_18), .B(n47), .C(Thlen_2), .D(n45), .Q(n207) );
  NAND41 U144 ( .A(n201), .B(n202), .C(n203), .D(n204), .Q(DAT_O_19) );
  NAND22 U145 ( .A(ctrl_19), .B(n38), .Q(n201) );
  AOI221 U146 ( .A(CBAR_19), .B(n2), .C(VBARb_19), .D(n49), .Q(n204) );
  AOI221 U147 ( .A(VBARa_19), .B(n47), .C(Thlen_3), .D(n45), .Q(n203) );
  NAND41 U148 ( .A(n193), .B(n194), .C(n195), .D(n196), .Q(DAT_O_20) );
  NAND22 U149 ( .A(ctrl_20), .B(n38), .Q(n193) );
  AOI221 U150 ( .A(CBAR_20), .B(n108), .C(VBARb_20), .D(n49), .Q(n196) );
  AOI221 U151 ( .A(VBARa_20), .B(n47), .C(Thlen_4), .D(n46), .Q(n195) );
  NAND41 U152 ( .A(n189), .B(n190), .C(n191), .D(n192), .Q(DAT_O_21) );
  NAND22 U153 ( .A(ctrl_21), .B(n38), .Q(n189) );
  AOI221 U154 ( .A(CBAR_21), .B(n2), .C(VBARb_21), .D(n50), .Q(n192) );
  AOI221 U155 ( .A(VBARa_21), .B(n47), .C(Thlen_5), .D(n46), .Q(n191) );
  NAND41 U156 ( .A(n185), .B(n186), .C(n187), .D(n188), .Q(DAT_O_22) );
  NAND22 U157 ( .A(ctrl_22), .B(n38), .Q(n185) );
  AOI221 U158 ( .A(CBAR_22), .B(n2), .C(VBARb_22), .D(n50), .Q(n188) );
  AOI221 U159 ( .A(VBARa_22), .B(n47), .C(Thlen_6), .D(n46), .Q(n187) );
  NAND41 U160 ( .A(n181), .B(n182), .C(n183), .D(n184), .Q(DAT_O_23) );
  NAND22 U161 ( .A(ctrl_23), .B(n38), .Q(n181) );
  AOI221 U162 ( .A(CBAR_23), .B(n2), .C(VBARb_23), .D(n50), .Q(n184) );
  AOI221 U163 ( .A(VBARa_23), .B(n47), .C(Thlen_7), .D(n46), .Q(n183) );
  NAND41 U164 ( .A(n177), .B(n178), .C(n179), .D(n180), .Q(DAT_O_24) );
  NAND22 U165 ( .A(ctrl_24), .B(n38), .Q(n177) );
  AOI221 U166 ( .A(CBAR_24), .B(n2), .C(VBARb_24), .D(n50), .Q(n180) );
  AOI221 U167 ( .A(VBARa_24), .B(n47), .C(Thlen_8), .D(n46), .Q(n179) );
  NAND41 U168 ( .A(n173), .B(n174), .C(n175), .D(n176), .Q(DAT_O_25) );
  NAND22 U169 ( .A(ctrl_25), .B(n38), .Q(n173) );
  AOI221 U170 ( .A(CBAR_25), .B(n108), .C(VBARb_25), .D(n50), .Q(n176) );
  AOI221 U171 ( .A(VBARa_25), .B(n47), .C(Thlen_9), .D(n46), .Q(n175) );
  NAND41 U172 ( .A(n169), .B(n170), .C(n171), .D(n172), .Q(DAT_O_26) );
  NAND22 U173 ( .A(ctrl_26), .B(n38), .Q(n169) );
  AOI221 U174 ( .A(CBAR_26), .B(n2), .C(VBARb_26), .D(n50), .Q(n172) );
  AOI221 U175 ( .A(VBARa_26), .B(n47), .C(Thlen_10), .D(n46), .Q(n171) );
  NAND41 U176 ( .A(n165), .B(n166), .C(n167), .D(n168), .Q(DAT_O_27) );
  NAND22 U177 ( .A(ctrl_27), .B(n37), .Q(n165) );
  AOI221 U178 ( .A(CBAR_27), .B(n108), .C(VBARb_27), .D(n50), .Q(n168) );
  AOI221 U179 ( .A(VBARa_27), .B(n48), .C(Thlen_11), .D(n45), .Q(n167) );
  NAND41 U180 ( .A(n161), .B(n162), .C(n163), .D(n164), .Q(DAT_O_28) );
  NAND22 U181 ( .A(ctrl_28), .B(n37), .Q(n161) );
  AOI221 U182 ( .A(CBAR_28), .B(n2), .C(VBARb_28), .D(n50), .Q(n164) );
  AOI221 U183 ( .A(VBARa_28), .B(n48), .C(Thlen_12), .D(n100), .Q(n163) );
  NAND41 U184 ( .A(n157), .B(n158), .C(n159), .D(n160), .Q(DAT_O_29) );
  NAND22 U185 ( .A(ctrl_29), .B(n37), .Q(n157) );
  AOI221 U186 ( .A(CBAR_29), .B(n2), .C(VBARb_29), .D(n49), .Q(n160) );
  AOI221 U187 ( .A(VBARa_29), .B(n48), .C(Thlen_13), .D(n100), .Q(n159) );
  NAND41 U188 ( .A(n149), .B(n150), .C(n151), .D(n152), .Q(DAT_O_30) );
  NAND22 U189 ( .A(ctrl_30), .B(n37), .Q(n149) );
  AOI221 U190 ( .A(CBAR_30), .B(n2), .C(VBARb_30), .D(n94), .Q(n152) );
  AOI221 U191 ( .A(VBARa_30), .B(n48), .C(Thlen_14), .D(n100), .Q(n151) );
  NAND41 U192 ( .A(n145), .B(n146), .C(n147), .D(n148), .Q(DAT_O_31) );
  NAND22 U193 ( .A(ctrl_31), .B(n37), .Q(n145) );
  AOI221 U194 ( .A(CBAR_31), .B(n2), .C(VBARb_31), .D(n94), .Q(n148) );
  AOI221 U195 ( .A(VBARa_31), .B(n48), .C(Thlen_15), .D(n100), .Q(n147) );
  NAND41 U196 ( .A(n197), .B(n198), .C(n199), .D(n200), .Q(DAT_O_2) );
  NAND22 U197 ( .A(ctrl_2_1), .B(n38), .Q(n198) );
  AOI221 U198 ( .A(VBARb_2), .B(n49), .C(VBARa_2), .D(n48), .Q(n200) );
  AOI221 U199 ( .A(Tvlen_2), .B(n45), .C(Tvgate_2), .D(n43), .Q(n199) );
  NAND41 U200 ( .A(n153), .B(n154), .C(n155), .D(n156), .Q(DAT_O_3) );
  NAND22 U201 ( .A(ctrl_3_1), .B(n37), .Q(n154) );
  AOI221 U202 ( .A(VBARb_3), .B(n49), .C(VBARa_3), .D(n48), .Q(n156) );
  AOI221 U203 ( .A(Tvlen_3), .B(n45), .C(Tvgate_3), .D(n43), .Q(n155) );
  NAND41 U204 ( .A(n129), .B(n130), .C(n131), .D(n132), .Q(DAT_O_7) );
  NAND22 U205 ( .A(VBL_0), .B(n37), .Q(n130) );
  AOI221 U206 ( .A(VBARb_7), .B(n50), .C(VBARa_7), .D(n96), .Q(n132) );
  AOI221 U207 ( .A(Tvlen_7), .B(n46), .C(Tvgate_7), .D(n43), .Q(n131) );
  NAND41 U208 ( .A(n125), .B(n126), .C(n127), .D(n128), .Q(DAT_O_8) );
  NAND22 U209 ( .A(VBL_1), .B(n37), .Q(n126) );
  AOI221 U210 ( .A(VBARb_8), .B(n50), .C(VBARa_8), .D(n96), .Q(n128) );
  AOI221 U211 ( .A(Tvlen_8), .B(n46), .C(Tvgate_8), .D(n43), .Q(n127) );
  NAND41 U212 ( .A(n120), .B(n121), .C(n122), .D(n123), .Q(DAT_O_9) );
  NAND22 U213 ( .A(CD_0), .B(n37), .Q(n121) );
  AOI221 U214 ( .A(VBARb_9), .B(n50), .C(VBARa_9), .D(n96), .Q(n123) );
  AOI221 U215 ( .A(Tvlen_9), .B(n46), .C(Tvgate_9), .D(n43), .Q(n122) );
  INV3 U216 ( .A(n63), .Q(n310) );
  AOI211 U217 ( .A(n320), .B(n50), .C(RST_I), .Q(n63) );
  INV3 U218 ( .A(n95), .Q(n309) );
  AOI211 U219 ( .A(n320), .B(n48), .C(RST_I), .Q(n95) );
  INV3 U220 ( .A(n101), .Q(n307) );
  AOI211 U221 ( .A(n320), .B(n44), .C(RST_I), .Q(n101) );
  INV3 U222 ( .A(n105), .Q(n305) );
  AOI211 U223 ( .A(n320), .B(n39), .C(RST_I), .Q(n105) );
  INV3 U224 ( .A(n103), .Q(n306) );
  AOI211 U225 ( .A(n320), .B(n41), .C(RST_I), .Q(n103) );
  OAI2111 U226 ( .A(n42), .B(n34), .C(n243), .D(n244), .Q(DAT_O_0) );
  AOI221 U227 ( .A(Tvlen_0), .B(n46), .C(Tvgate_0), .D(n43), .Q(n243) );
  AOI221 U228 ( .A(n124), .B(stat_0), .C(Ven), .D(n39), .Q(n244) );
  OAI2111 U229 ( .A(n42), .B(n33), .C(n241), .D(n242), .Q(DAT_O_1) );
  AOI221 U230 ( .A(Tvlen_1), .B(n45), .C(Tvgate_1), .D(n43), .Q(n241) );
  AOI221 U231 ( .A(n124), .B(stat_1), .C(ctrl_1_1), .D(n39), .Q(n242) );
  AOI221 U232 ( .A(stat_16), .B(n124), .C(ctrl_16), .D(n39), .Q(n213) );
  INV3 U233 ( .A(n107), .Q(n304) );
  AOI211 U234 ( .A(n320), .B(n108), .C(RST_I), .Q(n107) );
  INV3 U235 ( .A(ADR_I_3), .Q(n312) );
  INV3 U236 ( .A(ADR_I_4), .Q(n311) );
  INV3 U237 ( .A(ADR_I_2), .Q(n313) );
  AOI221 U238 ( .A(Thgate_4), .B(n41), .C(n124), .D(stat_4), .Q(n141) );
  AOI221 U239 ( .A(Thgate_5), .B(n41), .C(n124), .D(stat_5), .Q(n137) );
  AOI221 U240 ( .A(Thgate_6), .B(n41), .C(n124), .D(stat_6), .Q(n133) );
  AOI221 U241 ( .A(Tvgate_10), .B(n43), .C(Thgate_10), .D(n40), .Q(n238) );
  AOI221 U242 ( .A(Tvsync_5), .B(n43), .C(Thsync_5), .D(n41), .Q(n158) );
  AOI221 U243 ( .A(Tvsync_7), .B(n43), .C(Thsync_7), .D(n41), .Q(n146) );
  AOI221 U244 ( .A(Tvgdel_1), .B(n44), .C(Thgdel_1), .D(n40), .Q(n210) );
  AOI221 U245 ( .A(Tvgdel_2), .B(n44), .C(Thgdel_2), .D(n40), .Q(n206) );
  AOI221 U246 ( .A(Tvgdel_3), .B(n44), .C(Thgdel_3), .D(n40), .Q(n202) );
  AOI221 U247 ( .A(Tvgdel_4), .B(n44), .C(Thgdel_4), .D(n41), .Q(n194) );
  AOI221 U248 ( .A(Tvgdel_5), .B(n44), .C(Thgdel_5), .D(n41), .Q(n190) );
  AOI221 U249 ( .A(Tvgdel_6), .B(n44), .C(Thgdel_6), .D(n41), .Q(n186) );
  AOI221 U250 ( .A(Tvgdel_7), .B(n43), .C(Thgdel_7), .D(n41), .Q(n182) );
  AOI221 U251 ( .A(Tvsync_0), .B(n44), .C(Thsync_0), .D(n41), .Q(n178) );
  AOI221 U252 ( .A(Tvsync_1), .B(n102), .C(Thsync_1), .D(n41), .Q(n174) );
  AOI221 U253 ( .A(Tvsync_2), .B(n102), .C(Thsync_2), .D(n41), .Q(n170) );
  AOI221 U254 ( .A(Tvsync_3), .B(n102), .C(Thsync_3), .D(n41), .Q(n166) );
  AOI221 U255 ( .A(Tvsync_4), .B(n102), .C(Thsync_4), .D(n41), .Q(n162) );
  AOI221 U256 ( .A(Tvsync_6), .B(n102), .C(Thsync_6), .D(n41), .Q(n150) );
  AOI221 U257 ( .A(Tvgate_11), .B(n44), .C(Thgate_11), .D(n40), .Q(n234) );
  AOI221 U258 ( .A(Tvgate_12), .B(n44), .C(Thgate_12), .D(n40), .Q(n230) );
  AOI221 U259 ( .A(Tvgate_13), .B(n44), .C(Thgate_13), .D(n40), .Q(n226) );
  AOI221 U260 ( .A(Tvgate_14), .B(n44), .C(Thgate_14), .D(n40), .Q(n222) );
  AOI221 U261 ( .A(Tvgate_15), .B(n44), .C(Thgate_15), .D(n40), .Q(n218) );
  INV3 U262 ( .A(n97), .Q(n308) );
  AOI211 U263 ( .A(n320), .B(n46), .C(RST_I), .Q(n97) );
  INV3 U264 ( .A(n104), .Q(n42) );
  NOR31 U265 ( .A(ADR_I_2), .B(ADR_I_4), .C(n312), .Q(n104) );
  NAND22 U266 ( .A(Thgate_2), .B(n40), .Q(n197) );
  NAND22 U267 ( .A(Thgate_3), .B(n40), .Q(n153) );
  NAND22 U268 ( .A(Thgate_7), .B(n40), .Q(n129) );
  NAND22 U269 ( .A(Thgate_8), .B(n40), .Q(n125) );
  NAND22 U270 ( .A(Thgate_9), .B(n40), .Q(n120) );
  INV3 U271 ( .A(CYC_I), .Q(n322) );
  INV3 U272 ( .A(STB_I), .Q(n321) );
  AOI211 U273 ( .A(n270), .B(n116), .C(RST_I), .Q(N66) );
  INV3 U274 ( .A(sint_in), .Q(n270) );
  INV3 U275 ( .A(DAT_I_0), .Q(n318) );
  AOI211 U276 ( .A(n323), .B(n115), .C(RST_I), .Q(N67) );
  INV3 U277 ( .A(luint_in), .Q(n323) );
  INV3 U278 ( .A(DAT_I_1), .Q(n317) );
  AOI211 U279 ( .A(n266), .B(n114), .C(RST_I), .Q(N68) );
  INV3 U280 ( .A(vint_in), .Q(n266) );
  INV3 U281 ( .A(DAT_I_4), .Q(n316) );
  AOI211 U282 ( .A(n265), .B(n113), .C(RST_I), .Q(N69) );
  INV3 U283 ( .A(hint_in), .Q(n265) );
  INV3 U284 ( .A(DAT_I_5), .Q(n315) );
  AOI211 U285 ( .A(n267), .B(n112), .C(RST_I), .Q(N70) );
  INV3 U286 ( .A(bsint_in), .Q(n267) );
  INV3 U287 ( .A(DAT_I_6), .Q(n314) );
  NAND22 U288 ( .A(n117), .B(n118), .Q(INTA_O) );
  AOI221 U289 ( .A(stat_5), .B(ctrl_2_1), .C(stat_6), .D(ctrl_3_1), .Q(n117)
         );
  AOI2111 U290 ( .A(stat_4), .B(ctrl_1_1), .C(stat_1), .D(stat_0), .Q(n118) );
  INV3 U291 ( .A(n88), .Q(n297) );
  NAND22 U292 ( .A(DAT_I_26), .B(n4), .Q(n88) );
  INV3 U293 ( .A(n89), .Q(n298) );
  NAND22 U294 ( .A(DAT_I_27), .B(n4), .Q(n89) );
  INV3 U295 ( .A(n90), .Q(n299) );
  NAND22 U296 ( .A(DAT_I_28), .B(n4), .Q(n90) );
  INV3 U297 ( .A(n91), .Q(n300) );
  NAND22 U298 ( .A(DAT_I_29), .B(n4), .Q(n91) );
  INV3 U299 ( .A(n92), .Q(n301) );
  NAND22 U300 ( .A(DAT_I_30), .B(n4), .Q(n92) );
  INV3 U301 ( .A(n93), .Q(n302) );
  NAND22 U302 ( .A(DAT_I_31), .B(n4), .Q(n93) );
  INV3 U303 ( .A(n64), .Q(n273) );
  NAND22 U304 ( .A(DAT_I_2), .B(n3), .Q(n64) );
  INV3 U305 ( .A(n65), .Q(n274) );
  NAND22 U306 ( .A(DAT_I_3), .B(n3), .Q(n65) );
  INV3 U307 ( .A(n66), .Q(n275) );
  NAND22 U308 ( .A(DAT_I_4), .B(n3), .Q(n66) );
  INV3 U309 ( .A(n67), .Q(n276) );
  NAND22 U310 ( .A(DAT_I_5), .B(n3), .Q(n67) );
  INV3 U311 ( .A(n68), .Q(n277) );
  NAND22 U312 ( .A(DAT_I_6), .B(n3), .Q(n68) );
  INV3 U313 ( .A(n69), .Q(n278) );
  NAND22 U314 ( .A(DAT_I_7), .B(n3), .Q(n69) );
  INV3 U315 ( .A(n70), .Q(n279) );
  NAND22 U316 ( .A(DAT_I_8), .B(n3), .Q(n70) );
  INV3 U317 ( .A(n71), .Q(n280) );
  NAND22 U318 ( .A(DAT_I_9), .B(n3), .Q(n71) );
  INV3 U319 ( .A(n72), .Q(n281) );
  NAND22 U320 ( .A(DAT_I_10), .B(n3), .Q(n72) );
  INV3 U321 ( .A(RST_I), .Q(n303) );
  INV3 U322 ( .A(n98), .Q(n271) );
  NAND22 U323 ( .A(DAT_I_0), .B(n3), .Q(n98) );
  INV3 U324 ( .A(n99), .Q(n272) );
  NAND22 U325 ( .A(DAT_I_1), .B(n3), .Q(n99) );
  INV3 U326 ( .A(n73), .Q(n282) );
  NAND22 U327 ( .A(DAT_I_11), .B(n3), .Q(n73) );
  INV3 U328 ( .A(n74), .Q(n283) );
  NAND22 U329 ( .A(DAT_I_12), .B(n3), .Q(n74) );
  INV3 U330 ( .A(n75), .Q(n284) );
  NAND22 U331 ( .A(DAT_I_13), .B(n4), .Q(n75) );
  INV3 U332 ( .A(n76), .Q(n285) );
  NAND22 U333 ( .A(DAT_I_14), .B(n4), .Q(n76) );
  INV3 U334 ( .A(n77), .Q(n286) );
  NAND22 U335 ( .A(DAT_I_15), .B(n4), .Q(n77) );
  INV3 U336 ( .A(n78), .Q(n287) );
  NAND22 U337 ( .A(DAT_I_16), .B(n4), .Q(n78) );
  INV3 U338 ( .A(n79), .Q(n288) );
  NAND22 U339 ( .A(DAT_I_17), .B(n4), .Q(n79) );
  INV3 U340 ( .A(n80), .Q(n289) );
  NAND22 U341 ( .A(DAT_I_18), .B(n303), .Q(n80) );
  INV3 U342 ( .A(n81), .Q(n290) );
  NAND22 U343 ( .A(DAT_I_19), .B(n303), .Q(n81) );
  INV3 U344 ( .A(n82), .Q(n291) );
  NAND22 U345 ( .A(DAT_I_20), .B(n303), .Q(n82) );
  INV3 U346 ( .A(n83), .Q(n292) );
  NAND22 U347 ( .A(DAT_I_21), .B(n303), .Q(n83) );
  INV3 U348 ( .A(n84), .Q(n293) );
  NAND22 U349 ( .A(DAT_I_22), .B(n303), .Q(n84) );
  INV3 U350 ( .A(n85), .Q(n294) );
  NAND22 U351 ( .A(DAT_I_23), .B(n303), .Q(n85) );
  INV3 U352 ( .A(n86), .Q(n295) );
  NAND22 U353 ( .A(DAT_I_24), .B(n303), .Q(n86) );
  INV3 U354 ( .A(n87), .Q(n296) );
  NAND22 U355 ( .A(DAT_I_25), .B(n303), .Q(n87) );
  INV3 U356 ( .A(n111), .Q(n269) );
  NAND22 U357 ( .A(n4), .B(AVMP), .Q(n111) );
  INV3 U358 ( .A(n110), .Q(n268) );
  NAND22 U359 ( .A(n4), .B(ACMP), .Q(n110) );
  BUF2 U360 ( .A(NRESET), .Q(n58) );
  BUF2 U361 ( .A(NRESET), .Q(n59) );
  BUF2 U362 ( .A(NRESET), .Q(n61) );
  BUF2 U363 ( .A(NRESET), .Q(n60) );
endmodule


module Tgen ( clk, rst, HSyncL, .Thsync({Thsync_7, Thsync_6, Thsync_5, 
        Thsync_4, Thsync_3, Thsync_2, Thsync_1, Thsync_0}), .Thgdel({Thgdel_7, 
        Thgdel_6, Thgdel_5, Thgdel_4, Thgdel_3, Thgdel_2, Thgdel_1, Thgdel_0}), 
    .Thgate({Thgate_15, Thgate_14, Thgate_13, Thgate_12, Thgate_11, Thgate_10, 
        Thgate_9, Thgate_8, Thgate_7, Thgate_6, Thgate_5, Thgate_4, Thgate_3, 
        Thgate_2, Thgate_1, Thgate_0}), .Thlen({Thlen_15, Thlen_14, Thlen_13, 
        Thlen_12, Thlen_11, Thlen_10, Thlen_9, Thlen_8, Thlen_7, Thlen_6, 
        Thlen_5, Thlen_4, Thlen_3, Thlen_2, Thlen_1, Thlen_0}), VSyncL, 
    .Tvsync({Tvsync_7, Tvsync_6, Tvsync_5, Tvsync_4, Tvsync_3, Tvsync_2, 
        Tvsync_1, Tvsync_0}), .Tvgdel({Tvgdel_7, Tvgdel_6, Tvgdel_5, Tvgdel_4, 
        Tvgdel_3, Tvgdel_2, Tvgdel_1, Tvgdel_0}), .Tvgate({Tvgate_15, 
        Tvgate_14, Tvgate_13, Tvgate_12, Tvgate_11, Tvgate_10, Tvgate_9, 
        Tvgate_8, Tvgate_7, Tvgate_6, Tvgate_5, Tvgate_4, Tvgate_3, Tvgate_2, 
        Tvgate_1, Tvgate_0}), .Tvlen({Tvlen_15, Tvlen_14, Tvlen_13, Tvlen_12, 
        Tvlen_11, Tvlen_10, Tvlen_9, Tvlen_8, Tvlen_7, Tvlen_6, Tvlen_5, 
        Tvlen_4, Tvlen_3, Tvlen_2, Tvlen_1, Tvlen_0}), CSyncL, BlankL, eol, 
        eof, gate, Hsync, Vsync, Csync, Blank );
  input clk, rst, HSyncL, Thsync_7, Thsync_6, Thsync_5, Thsync_4, Thsync_3,
         Thsync_2, Thsync_1, Thsync_0, Thgdel_7, Thgdel_6, Thgdel_5, Thgdel_4,
         Thgdel_3, Thgdel_2, Thgdel_1, Thgdel_0, Thgate_15, Thgate_14,
         Thgate_13, Thgate_12, Thgate_11, Thgate_10, Thgate_9, Thgate_8,
         Thgate_7, Thgate_6, Thgate_5, Thgate_4, Thgate_3, Thgate_2, Thgate_1,
         Thgate_0, Thlen_15, Thlen_14, Thlen_13, Thlen_12, Thlen_11, Thlen_10,
         Thlen_9, Thlen_8, Thlen_7, Thlen_6, Thlen_5, Thlen_4, Thlen_3,
         Thlen_2, Thlen_1, Thlen_0, VSyncL, Tvsync_7, Tvsync_6, Tvsync_5,
         Tvsync_4, Tvsync_3, Tvsync_2, Tvsync_1, Tvsync_0, Tvgdel_7, Tvgdel_6,
         Tvgdel_5, Tvgdel_4, Tvgdel_3, Tvgdel_2, Tvgdel_1, Tvgdel_0, Tvgate_15,
         Tvgate_14, Tvgate_13, Tvgate_12, Tvgate_11, Tvgate_10, Tvgate_9,
         Tvgate_8, Tvgate_7, Tvgate_6, Tvgate_5, Tvgate_4, Tvgate_3, Tvgate_2,
         Tvgate_1, Tvgate_0, Tvlen_15, Tvlen_14, Tvlen_13, Tvlen_12, Tvlen_11,
         Tvlen_10, Tvlen_9, Tvlen_8, Tvlen_7, Tvlen_6, Tvlen_5, Tvlen_4,
         Tvlen_3, Tvlen_2, Tvlen_1, Tvlen_0, CSyncL, BlankL;
  output eol, eof, gate, Hsync, Vsync, Csync, Blank;
  wire   iHsync, Hgate, iVsync, Vgate, n2, n3, n1;

  vtim hor_gen ( .clk(clk), .ena(n1), .rst(rst), .Tsync({Thsync_7, Thsync_6, 
        Thsync_5, Thsync_4, Thsync_3, Thsync_2, Thsync_1, Thsync_0}), .Tgdel({
        Thgdel_7, Thgdel_6, Thgdel_5, Thgdel_4, Thgdel_3, Thgdel_2, Thgdel_1, 
        Thgdel_0}), .Tgate({Thgate_15, Thgate_14, Thgate_13, Thgate_12, 
        Thgate_11, Thgate_10, Thgate_9, Thgate_8, Thgate_7, Thgate_6, Thgate_5, 
        Thgate_4, Thgate_3, Thgate_2, Thgate_1, Thgate_0}), .Tlen({Thlen_15, 
        Thlen_14, Thlen_13, Thlen_12, Thlen_11, Thlen_10, Thlen_9, Thlen_8, 
        Thlen_7, Thlen_6, Thlen_5, Thlen_4, Thlen_3, Thlen_2, Thlen_1, Thlen_0}), .Sync(iHsync), .Gate(Hgate), .Done(eol) );
  vtim ver_gen ( .clk(clk), .ena(eol), .rst(rst), .Tsync({Tvsync_7, Tvsync_6, 
        Tvsync_5, Tvsync_4, Tvsync_3, Tvsync_2, Tvsync_1, Tvsync_0}), .Tgdel({
        Tvgdel_7, Tvgdel_6, Tvgdel_5, Tvgdel_4, Tvgdel_3, Tvgdel_2, Tvgdel_1, 
        Tvgdel_0}), .Tgate({Tvgate_15, Tvgate_14, Tvgate_13, Tvgate_12, 
        Tvgate_11, Tvgate_10, Tvgate_9, Tvgate_8, Tvgate_7, Tvgate_6, Tvgate_5, 
        Tvgate_4, Tvgate_3, Tvgate_2, Tvgate_1, Tvgate_0}), .Tlen({Tvlen_15, 
        Tvlen_14, Tvlen_13, Tvlen_12, Tvlen_11, Tvlen_10, Tvlen_9, Tvlen_8, 
        Tvlen_7, Tvlen_6, Tvlen_5, Tvlen_4, Tvlen_3, Tvlen_2, Tvlen_1, Tvlen_0}), .Sync(iVsync), .Gate(Vgate), .Done(eof) );
  INV3 U2 ( .A(n2), .Q(gate) );
  NAND22 U3 ( .A(Vgate), .B(Hgate), .Q(n2) );
  XOR21 U4 ( .A(iHsync), .B(HSyncL), .Q(Hsync) );
  XOR21 U5 ( .A(iVsync), .B(VSyncL), .Q(Vsync) );
  XNR21 U6 ( .A(BlankL), .B(gate), .Q(Blank) );
  XNR21 U7 ( .A(CSyncL), .B(n3), .Q(Csync) );
  NOR21 U8 ( .A(iHsync), .B(iVsync), .Q(n3) );
  LOGIC1 U9 ( .Q(n1) );
endmodule


module Pgen ( mclk, pclk, ctrl_Ven, ctrl_HSyncL, .Thsync({Thsync_7, Thsync_6, 
        Thsync_5, Thsync_4, Thsync_3, Thsync_2, Thsync_1, Thsync_0}), 
    .Thgdel({Thgdel_7, Thgdel_6, Thgdel_5, Thgdel_4, Thgdel_3, Thgdel_2, 
        Thgdel_1, Thgdel_0}), .Thgate({Thgate_15, Thgate_14, Thgate_13, 
        Thgate_12, Thgate_11, Thgate_10, Thgate_9, Thgate_8, Thgate_7, 
        Thgate_6, Thgate_5, Thgate_4, Thgate_3, Thgate_2, Thgate_1, Thgate_0}), 
    .Thlen({Thlen_15, Thlen_14, Thlen_13, Thlen_12, Thlen_11, Thlen_10, 
        Thlen_9, Thlen_8, Thlen_7, Thlen_6, Thlen_5, Thlen_4, Thlen_3, Thlen_2, 
        Thlen_1, Thlen_0}), ctrl_VSyncL, .Tvsync({Tvsync_7, Tvsync_6, Tvsync_5, 
        Tvsync_4, Tvsync_3, Tvsync_2, Tvsync_1, Tvsync_0}), .Tvgdel({Tvgdel_7, 
        Tvgdel_6, Tvgdel_5, Tvgdel_4, Tvgdel_3, Tvgdel_2, Tvgdel_1, Tvgdel_0}), 
    .Tvgate({Tvgate_15, Tvgate_14, Tvgate_13, Tvgate_12, Tvgate_11, Tvgate_10, 
        Tvgate_9, Tvgate_8, Tvgate_7, Tvgate_6, Tvgate_5, Tvgate_4, Tvgate_3, 
        Tvgate_2, Tvgate_1, Tvgate_0}), .Tvlen({Tvlen_15, Tvlen_14, Tvlen_13, 
        Tvlen_12, Tvlen_11, Tvlen_10, Tvlen_9, Tvlen_8, Tvlen_7, Tvlen_6, 
        Tvlen_5, Tvlen_4, Tvlen_3, Tvlen_2, Tvlen_1, Tvlen_0}), ctrl_CSyncL, 
        ctrl_BlankL, eoh, eov, Gate, Hsync, Vsync, Csync, Blank );
  input mclk, pclk, ctrl_Ven, ctrl_HSyncL, Thsync_7, Thsync_6, Thsync_5,
         Thsync_4, Thsync_3, Thsync_2, Thsync_1, Thsync_0, Thgdel_7, Thgdel_6,
         Thgdel_5, Thgdel_4, Thgdel_3, Thgdel_2, Thgdel_1, Thgdel_0, Thgate_15,
         Thgate_14, Thgate_13, Thgate_12, Thgate_11, Thgate_10, Thgate_9,
         Thgate_8, Thgate_7, Thgate_6, Thgate_5, Thgate_4, Thgate_3, Thgate_2,
         Thgate_1, Thgate_0, Thlen_15, Thlen_14, Thlen_13, Thlen_12, Thlen_11,
         Thlen_10, Thlen_9, Thlen_8, Thlen_7, Thlen_6, Thlen_5, Thlen_4,
         Thlen_3, Thlen_2, Thlen_1, Thlen_0, ctrl_VSyncL, Tvsync_7, Tvsync_6,
         Tvsync_5, Tvsync_4, Tvsync_3, Tvsync_2, Tvsync_1, Tvsync_0, Tvgdel_7,
         Tvgdel_6, Tvgdel_5, Tvgdel_4, Tvgdel_3, Tvgdel_2, Tvgdel_1, Tvgdel_0,
         Tvgate_15, Tvgate_14, Tvgate_13, Tvgate_12, Tvgate_11, Tvgate_10,
         Tvgate_9, Tvgate_8, Tvgate_7, Tvgate_6, Tvgate_5, Tvgate_4, Tvgate_3,
         Tvgate_2, Tvgate_1, Tvgate_0, Tvlen_15, Tvlen_14, Tvlen_13, Tvlen_12,
         Tvlen_11, Tvlen_10, Tvlen_9, Tvlen_8, Tvlen_7, Tvlen_6, Tvlen_5,
         Tvlen_4, Tvlen_3, Tvlen_2, Tvlen_1, Tvlen_0, ctrl_CSyncL, ctrl_BlankL;
  output eoh, eov, Gate, Hsync, Vsync, Csync, Blank;
  wire   nVen, eol, eof, seol, dseol, seof, dseof, N1, N2, n1, n2, n3;

  DF3 nVen_reg ( .D(n3), .C(pclk), .Q(nVen) );
  DF3 seol_reg ( .D(eol), .C(mclk), .Q(seol), .QN(n1) );
  DF3 dseol_reg ( .D(seol), .C(mclk), .Q(dseol) );
  DF3 seof_reg ( .D(eof), .C(mclk), .Q(seof), .QN(n2) );
  DF3 dseof_reg ( .D(seof), .C(mclk), .Q(dseof) );
  DF3 eoh_reg ( .D(N1), .C(mclk), .Q(eoh) );
  DF3 eov_reg ( .D(N2), .C(mclk), .Q(eov) );
  Tgen vtgen ( .clk(pclk), .rst(nVen), .HSyncL(ctrl_HSyncL), .Thsync({Thsync_7, 
        Thsync_6, Thsync_5, Thsync_4, Thsync_3, Thsync_2, Thsync_1, Thsync_0}), 
        .Thgdel({Thgdel_7, Thgdel_6, Thgdel_5, Thgdel_4, Thgdel_3, Thgdel_2, 
        Thgdel_1, Thgdel_0}), .Thgate({Thgate_15, Thgate_14, Thgate_13, 
        Thgate_12, Thgate_11, Thgate_10, Thgate_9, Thgate_8, Thgate_7, 
        Thgate_6, Thgate_5, Thgate_4, Thgate_3, Thgate_2, Thgate_1, Thgate_0}), 
        .Thlen({Thlen_15, Thlen_14, Thlen_13, Thlen_12, Thlen_11, Thlen_10, 
        Thlen_9, Thlen_8, Thlen_7, Thlen_6, Thlen_5, Thlen_4, Thlen_3, Thlen_2, 
        Thlen_1, Thlen_0}), .VSyncL(ctrl_VSyncL), .Tvsync({Tvsync_7, Tvsync_6, 
        Tvsync_5, Tvsync_4, Tvsync_3, Tvsync_2, Tvsync_1, Tvsync_0}), .Tvgdel(
        {Tvgdel_7, Tvgdel_6, Tvgdel_5, Tvgdel_4, Tvgdel_3, Tvgdel_2, Tvgdel_1, 
        Tvgdel_0}), .Tvgate({Tvgate_15, Tvgate_14, Tvgate_13, Tvgate_12, 
        Tvgate_11, Tvgate_10, Tvgate_9, Tvgate_8, Tvgate_7, Tvgate_6, Tvgate_5, 
        Tvgate_4, Tvgate_3, Tvgate_2, Tvgate_1, Tvgate_0}), .Tvlen({Tvlen_15, 
        Tvlen_14, Tvlen_13, Tvlen_12, Tvlen_11, Tvlen_10, Tvlen_9, Tvlen_8, 
        Tvlen_7, Tvlen_6, Tvlen_5, Tvlen_4, Tvlen_3, Tvlen_2, Tvlen_1, Tvlen_0}), .CSyncL(ctrl_CSyncL), .BlankL(ctrl_BlankL), .eol(eol), .eof(eof), .gate(
        Gate), .Hsync(Hsync), .Vsync(Vsync), .Csync(Csync), .Blank(Blank) );
  INV3 U3 ( .A(ctrl_Ven), .Q(n3) );
  NOR21 U4 ( .A(dseof), .B(n2), .Q(N2) );
  NOR21 U5 ( .A(dseol), .B(n1), .Q(N1) );
endmodule


module dual_ported_memory_AWIDTH8_DWIDTH24 ( rclk, wclk, .D({D_23, D_22, D_21, 
        D_20, D_19, D_18, D_17, D_16, D_15, D_14, D_13, D_12, D_11, D_10, D_9, 
        D_8, D_7, D_6, D_5, D_4, D_3, D_2, D_1, D_0}), .waddr({waddr_7, 
        waddr_6, waddr_5, waddr_4, waddr_3, waddr_2, waddr_1, waddr_0}), wreq, 
    .Q({Q_23, Q_22, Q_21, Q_20, Q_19, Q_18, Q_17, Q_16, Q_15, Q_14, Q_13, Q_12, 
        Q_11, Q_10, Q_9, Q_8, Q_7, Q_6, Q_5, Q_4, Q_3, Q_2, Q_1, Q_0}), 
    .raddr({raddr_7, raddr_6, raddr_5, raddr_4, raddr_3, raddr_2, raddr_1, 
        raddr_0}) );
  input rclk, wclk, D_23, D_22, D_21, D_20, D_19, D_18, D_17, D_16, D_15, D_14,
         D_13, D_12, D_11, D_10, D_9, D_8, D_7, D_6, D_5, D_4, D_3, D_2, D_1,
         D_0, waddr_7, waddr_6, waddr_5, waddr_4, waddr_3, waddr_2, waddr_1,
         waddr_0, wreq, raddr_7, raddr_6, raddr_5, raddr_4, raddr_3, raddr_2,
         raddr_1, raddr_0;
  output Q_23, Q_22, Q_21, Q_20, Q_19, Q_18, Q_17, Q_16, Q_15, Q_14, Q_13,
         Q_12, Q_11, Q_10, Q_9, Q_8, Q_7, Q_6, Q_5, Q_4, Q_3, Q_2, Q_1, Q_0;
  wire   N791, N792, N793, N794, N795, N796, N797, N798, N799, N800, N801,
         N802, N803, N804, N805, N806, N807, N808, N809, N810, N811, N812,
         N813, N814, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351;

  OAI222 U311 ( .A(n2472), .B(n11091), .C(n2448), .D(n6512), .Q(n6510) );
  OAI222 U312 ( .A(n2424), .B(n11089), .C(n2400), .D(n6514), .Q(n6509) );
  OAI222 U313 ( .A(n2376), .B(n11087), .C(n2352), .D(n6516), .Q(n6508) );
  OAI222 U314 ( .A(n2328), .B(n11085), .C(n2304), .D(n6518), .Q(n6507) );
  OAI222 U316 ( .A(n2664), .B(n11083), .C(n2640), .D(n6524), .Q(n6522) );
  OAI222 U317 ( .A(n2616), .B(n11081), .C(n2592), .D(n6526), .Q(n6521) );
  OAI222 U318 ( .A(n2568), .B(n11079), .C(n2544), .D(n6528), .Q(n6520) );
  OAI222 U319 ( .A(n2520), .B(n11077), .C(n2496), .D(n6530), .Q(n6519) );
  OAI222 U321 ( .A(n2856), .B(n11075), .C(n2832), .D(n6536), .Q(n6534) );
  OAI222 U322 ( .A(n2808), .B(n11073), .C(n2784), .D(n6538), .Q(n6533) );
  OAI222 U323 ( .A(n2760), .B(n11071), .C(n2736), .D(n6540), .Q(n6532) );
  OAI222 U324 ( .A(n2712), .B(n11069), .C(n2688), .D(n6542), .Q(n6531) );
  OAI222 U326 ( .A(n3048), .B(n11067), .C(n3024), .D(n6548), .Q(n6546) );
  OAI222 U327 ( .A(n3000), .B(n11065), .C(n2976), .D(n6550), .Q(n6545) );
  OAI222 U328 ( .A(n2952), .B(n11063), .C(n2928), .D(n6552), .Q(n6544) );
  OAI222 U329 ( .A(n2904), .B(n11061), .C(n2880), .D(n6554), .Q(n6543) );
  OAI222 U332 ( .A(n1704), .B(n11059), .C(n1680), .D(n6564), .Q(n6562) );
  OAI222 U333 ( .A(n1656), .B(n11057), .C(n1632), .D(n6566), .Q(n6561) );
  OAI222 U334 ( .A(n1608), .B(n11055), .C(n1584), .D(n6568), .Q(n6560) );
  OAI222 U335 ( .A(n1560), .B(n11053), .C(n1536), .D(n6570), .Q(n6559) );
  OAI222 U337 ( .A(n1896), .B(n11051), .C(n1872), .D(n6576), .Q(n6574) );
  OAI222 U338 ( .A(n1848), .B(n11049), .C(n1824), .D(n6578), .Q(n6573) );
  OAI222 U339 ( .A(n1800), .B(n11047), .C(n1776), .D(n6580), .Q(n6572) );
  OAI222 U340 ( .A(n1752), .B(n11045), .C(n1728), .D(n6582), .Q(n6571) );
  OAI222 U342 ( .A(n2088), .B(n11043), .C(n2064), .D(n6588), .Q(n6586) );
  OAI222 U343 ( .A(n2040), .B(n11041), .C(n2016), .D(n6590), .Q(n6585) );
  OAI222 U344 ( .A(n1992), .B(n11039), .C(n1968), .D(n6592), .Q(n6584) );
  OAI222 U345 ( .A(n1944), .B(n11037), .C(n1920), .D(n6594), .Q(n6583) );
  OAI222 U347 ( .A(n2280), .B(n11035), .C(n2256), .D(n6600), .Q(n6598) );
  OAI222 U348 ( .A(n2232), .B(n11033), .C(n2208), .D(n6602), .Q(n6597) );
  OAI222 U349 ( .A(n2184), .B(n11031), .C(n2160), .D(n6604), .Q(n6596) );
  OAI222 U350 ( .A(n2136), .B(n11029), .C(n2112), .D(n6606), .Q(n6595) );
  OAI222 U353 ( .A(n936), .B(n11027), .C(n912), .D(n6616), .Q(n6614) );
  OAI222 U354 ( .A(n888), .B(n11025), .C(n864), .D(n6618), .Q(n6613) );
  OAI222 U355 ( .A(n840), .B(n11023), .C(n816), .D(n6620), .Q(n6612) );
  OAI222 U356 ( .A(n792), .B(n11021), .C(n768), .D(n6622), .Q(n6611) );
  OAI222 U358 ( .A(n1128), .B(n11019), .C(n1104), .D(n6628), .Q(n6626) );
  OAI222 U359 ( .A(n1080), .B(n11017), .C(n1056), .D(n6630), .Q(n6625) );
  OAI222 U360 ( .A(n1032), .B(n11015), .C(n1008), .D(n6632), .Q(n6624) );
  OAI222 U361 ( .A(n984), .B(n11013), .C(n960), .D(n6634), .Q(n6623) );
  OAI222 U363 ( .A(n1320), .B(n11011), .C(n1296), .D(n6640), .Q(n6638) );
  OAI222 U364 ( .A(n1272), .B(n11009), .C(n1248), .D(n6642), .Q(n6637) );
  OAI222 U365 ( .A(n1224), .B(n11007), .C(n1200), .D(n6644), .Q(n6636) );
  OAI222 U366 ( .A(n1176), .B(n11005), .C(n1152), .D(n6646), .Q(n6635) );
  OAI222 U368 ( .A(n1512), .B(n11003), .C(n1488), .D(n6652), .Q(n6650) );
  OAI222 U369 ( .A(n1464), .B(n11001), .C(n1440), .D(n6654), .Q(n6649) );
  OAI222 U370 ( .A(n1416), .B(n10999), .C(n1392), .D(n6656), .Q(n6648) );
  OAI222 U371 ( .A(n1368), .B(n10997), .C(n1344), .D(n6658), .Q(n6647) );
  OAI222 U374 ( .A(n168), .B(n10995), .C(n144), .D(n6668), .Q(n6666) );
  OAI222 U375 ( .A(n120), .B(n10993), .C(n96), .D(n6670), .Q(n6665) );
  OAI222 U376 ( .A(n72), .B(n10991), .C(n48), .D(n6672), .Q(n6664) );
  OAI222 U377 ( .A(n24), .B(n10989), .C(n6144), .D(n6674), .Q(n6663) );
  OAI222 U379 ( .A(n360), .B(n10987), .C(n336), .D(n6680), .Q(n6678) );
  OAI222 U380 ( .A(n312), .B(n10985), .C(n288), .D(n6682), .Q(n6677) );
  OAI222 U381 ( .A(n264), .B(n10983), .C(n240), .D(n6684), .Q(n6676) );
  OAI222 U382 ( .A(n216), .B(n10981), .C(n192), .D(n6686), .Q(n6675) );
  OAI222 U384 ( .A(n552), .B(n10979), .C(n528), .D(n6692), .Q(n6690) );
  OAI222 U385 ( .A(n504), .B(n10977), .C(n480), .D(n6694), .Q(n6689) );
  OAI222 U386 ( .A(n456), .B(n10975), .C(n432), .D(n6696), .Q(n6688) );
  OAI222 U387 ( .A(n408), .B(n10973), .C(n384), .D(n6698), .Q(n6687) );
  OAI222 U389 ( .A(n744), .B(n10971), .C(n720), .D(n6704), .Q(n6702) );
  OAI222 U390 ( .A(n696), .B(n10969), .C(n672), .D(n6706), .Q(n6701) );
  OAI222 U391 ( .A(n648), .B(n10967), .C(n624), .D(n6708), .Q(n6700) );
  OAI222 U392 ( .A(n600), .B(n10965), .C(n576), .D(n6710), .Q(n6699) );
  OAI222 U396 ( .A(n5544), .B(n10963), .C(n5520), .D(n6724), .Q(n6722) );
  OAI222 U397 ( .A(n5496), .B(n10961), .C(n5472), .D(n6726), .Q(n6721) );
  OAI222 U398 ( .A(n5448), .B(n10959), .C(n5424), .D(n6728), .Q(n6720) );
  OAI222 U399 ( .A(n5400), .B(n10957), .C(n5376), .D(n6730), .Q(n6719) );
  OAI222 U401 ( .A(n5736), .B(n10955), .C(n5712), .D(n6736), .Q(n6734) );
  OAI222 U402 ( .A(n5688), .B(n10953), .C(n5664), .D(n6738), .Q(n6733) );
  OAI222 U403 ( .A(n5640), .B(n10951), .C(n5616), .D(n6740), .Q(n6732) );
  OAI222 U404 ( .A(n5592), .B(n10949), .C(n5568), .D(n6742), .Q(n6731) );
  OAI222 U406 ( .A(n5928), .B(n10947), .C(n5904), .D(n6748), .Q(n6746) );
  OAI222 U407 ( .A(n5880), .B(n10945), .C(n5856), .D(n6750), .Q(n6745) );
  OAI222 U408 ( .A(n5832), .B(n10943), .C(n5808), .D(n6752), .Q(n6744) );
  OAI222 U409 ( .A(n5784), .B(n10941), .C(n5760), .D(n6754), .Q(n6743) );
  OAI222 U411 ( .A(n6120), .B(n10939), .C(n6096), .D(n6760), .Q(n6758) );
  OAI222 U412 ( .A(n6072), .B(n10937), .C(n6048), .D(n6762), .Q(n6757) );
  OAI222 U413 ( .A(n6024), .B(n10935), .C(n6000), .D(n6764), .Q(n6756) );
  OAI222 U414 ( .A(n5976), .B(n10933), .C(n5952), .D(n6766), .Q(n6755) );
  OAI222 U417 ( .A(n4776), .B(n10931), .C(n4752), .D(n6776), .Q(n6774) );
  OAI222 U418 ( .A(n4728), .B(n10929), .C(n4704), .D(n6778), .Q(n6773) );
  OAI222 U419 ( .A(n4680), .B(n10927), .C(n4656), .D(n6780), .Q(n6772) );
  OAI222 U420 ( .A(n4632), .B(n10925), .C(n4608), .D(n6782), .Q(n6771) );
  OAI222 U422 ( .A(n4968), .B(n10923), .C(n4944), .D(n6788), .Q(n6786) );
  OAI222 U423 ( .A(n4920), .B(n10921), .C(n4896), .D(n6790), .Q(n6785) );
  OAI222 U424 ( .A(n4872), .B(n10919), .C(n4848), .D(n6792), .Q(n6784) );
  OAI222 U425 ( .A(n4824), .B(n10917), .C(n4800), .D(n6794), .Q(n6783) );
  OAI222 U427 ( .A(n5160), .B(n10915), .C(n5136), .D(n6800), .Q(n6798) );
  OAI222 U428 ( .A(n5112), .B(n10913), .C(n5088), .D(n6802), .Q(n6797) );
  OAI222 U429 ( .A(n5064), .B(n10911), .C(n5040), .D(n6804), .Q(n6796) );
  OAI222 U430 ( .A(n5016), .B(n10909), .C(n4992), .D(n6806), .Q(n6795) );
  OAI222 U432 ( .A(n5352), .B(n10907), .C(n5328), .D(n6812), .Q(n6810) );
  OAI222 U433 ( .A(n5304), .B(n10905), .C(n5280), .D(n6814), .Q(n6809) );
  OAI222 U434 ( .A(n5256), .B(n10903), .C(n5232), .D(n6816), .Q(n6808) );
  OAI222 U435 ( .A(n5208), .B(n10901), .C(n5184), .D(n6818), .Q(n6807) );
  OAI222 U438 ( .A(n4008), .B(n10899), .C(n3984), .D(n6828), .Q(n6826) );
  OAI222 U439 ( .A(n3960), .B(n10897), .C(n3936), .D(n6830), .Q(n6825) );
  OAI222 U440 ( .A(n3912), .B(n10895), .C(n3888), .D(n6832), .Q(n6824) );
  OAI222 U441 ( .A(n3864), .B(n10893), .C(n3840), .D(n6834), .Q(n6823) );
  OAI222 U443 ( .A(n4200), .B(n10891), .C(n4176), .D(n6840), .Q(n6838) );
  OAI222 U444 ( .A(n4152), .B(n10889), .C(n4128), .D(n6842), .Q(n6837) );
  OAI222 U445 ( .A(n4104), .B(n10887), .C(n4080), .D(n6844), .Q(n6836) );
  OAI222 U446 ( .A(n4056), .B(n10885), .C(n4032), .D(n6846), .Q(n6835) );
  OAI222 U448 ( .A(n4392), .B(n10883), .C(n4368), .D(n6852), .Q(n6850) );
  OAI222 U449 ( .A(n4344), .B(n10881), .C(n4320), .D(n6854), .Q(n6849) );
  OAI222 U450 ( .A(n4296), .B(n6191), .C(n4272), .D(n6856), .Q(n6848) );
  OAI222 U451 ( .A(n4248), .B(n6189), .C(n4224), .D(n6858), .Q(n6847) );
  OAI222 U453 ( .A(n4584), .B(n6187), .C(n4560), .D(n6864), .Q(n6862) );
  OAI222 U454 ( .A(n4536), .B(n6185), .C(n4512), .D(n6866), .Q(n6861) );
  OAI222 U455 ( .A(n4488), .B(n6183), .C(n4464), .D(n6868), .Q(n6860) );
  OAI222 U456 ( .A(n4440), .B(n6181), .C(n4416), .D(n6870), .Q(n6859) );
  OAI222 U459 ( .A(n3240), .B(n6179), .C(n3216), .D(n6880), .Q(n6878) );
  OAI222 U460 ( .A(n3192), .B(n6177), .C(n3168), .D(n6882), .Q(n6877) );
  OAI222 U461 ( .A(n3144), .B(n6175), .C(n3120), .D(n6884), .Q(n6876) );
  OAI222 U462 ( .A(n3096), .B(n6173), .C(n3072), .D(n6886), .Q(n6875) );
  OAI222 U464 ( .A(n3432), .B(n6171), .C(n3408), .D(n6892), .Q(n6890) );
  OAI222 U465 ( .A(n3384), .B(n6169), .C(n3360), .D(n6894), .Q(n6889) );
  OAI222 U466 ( .A(n3336), .B(n6167), .C(n3312), .D(n6896), .Q(n6888) );
  OAI222 U467 ( .A(n3288), .B(n6165), .C(n3264), .D(n6898), .Q(n6887) );
  OAI222 U469 ( .A(n3624), .B(n6163), .C(n3600), .D(n6904), .Q(n6902) );
  OAI222 U470 ( .A(n3576), .B(n6161), .C(n3552), .D(n6906), .Q(n6901) );
  OAI222 U471 ( .A(n3528), .B(n6159), .C(n3504), .D(n6908), .Q(n6900) );
  OAI222 U472 ( .A(n3480), .B(n6157), .C(n3456), .D(n6910), .Q(n6899) );
  OAI222 U474 ( .A(n3816), .B(n6155), .C(n3792), .D(n6916), .Q(n6914) );
  OAI222 U475 ( .A(n3768), .B(n6153), .C(n3744), .D(n6918), .Q(n6913) );
  OAI222 U476 ( .A(n3720), .B(n6151), .C(n3696), .D(n6920), .Q(n6912) );
  OAI222 U477 ( .A(n3672), .B(n6149), .C(n3648), .D(n6922), .Q(n6911) );
  OAI222 U482 ( .A(n2471), .B(n11091), .C(n2447), .D(n6512), .Q(n6936) );
  OAI222 U483 ( .A(n2423), .B(n11089), .C(n2399), .D(n6514), .Q(n6935) );
  OAI222 U484 ( .A(n2375), .B(n11087), .C(n2351), .D(n6516), .Q(n6934) );
  OAI222 U485 ( .A(n2327), .B(n11085), .C(n2303), .D(n6518), .Q(n6933) );
  OAI222 U487 ( .A(n2663), .B(n11083), .C(n2639), .D(n6524), .Q(n6940) );
  OAI222 U488 ( .A(n2615), .B(n11081), .C(n2591), .D(n6526), .Q(n6939) );
  OAI222 U489 ( .A(n2567), .B(n11079), .C(n2543), .D(n6528), .Q(n6938) );
  OAI222 U490 ( .A(n2519), .B(n11077), .C(n2495), .D(n6530), .Q(n6937) );
  OAI222 U492 ( .A(n2855), .B(n11075), .C(n2831), .D(n6536), .Q(n6944) );
  OAI222 U493 ( .A(n2807), .B(n11073), .C(n2783), .D(n6538), .Q(n6943) );
  OAI222 U494 ( .A(n2759), .B(n11071), .C(n2735), .D(n6540), .Q(n6942) );
  OAI222 U495 ( .A(n2711), .B(n11069), .C(n2687), .D(n6542), .Q(n6941) );
  OAI222 U497 ( .A(n3047), .B(n11067), .C(n3023), .D(n6548), .Q(n6948) );
  OAI222 U498 ( .A(n2999), .B(n11065), .C(n2975), .D(n6550), .Q(n6947) );
  OAI222 U499 ( .A(n2951), .B(n11063), .C(n2927), .D(n6552), .Q(n6946) );
  OAI222 U500 ( .A(n2903), .B(n11061), .C(n2879), .D(n6554), .Q(n6945) );
  OAI222 U503 ( .A(n1703), .B(n11059), .C(n1679), .D(n6564), .Q(n6956) );
  OAI222 U504 ( .A(n1655), .B(n11057), .C(n1631), .D(n6566), .Q(n6955) );
  OAI222 U505 ( .A(n1607), .B(n11055), .C(n1583), .D(n6568), .Q(n6954) );
  OAI222 U506 ( .A(n1559), .B(n11053), .C(n1535), .D(n6570), .Q(n6953) );
  OAI222 U508 ( .A(n1895), .B(n11051), .C(n1871), .D(n6576), .Q(n6960) );
  OAI222 U509 ( .A(n1847), .B(n11049), .C(n1823), .D(n6578), .Q(n6959) );
  OAI222 U510 ( .A(n1799), .B(n11047), .C(n1775), .D(n6580), .Q(n6958) );
  OAI222 U511 ( .A(n1751), .B(n11045), .C(n1727), .D(n6582), .Q(n6957) );
  OAI222 U513 ( .A(n2087), .B(n11043), .C(n2063), .D(n6588), .Q(n6964) );
  OAI222 U514 ( .A(n2039), .B(n11041), .C(n2015), .D(n6590), .Q(n6963) );
  OAI222 U515 ( .A(n1991), .B(n11039), .C(n1967), .D(n6592), .Q(n6962) );
  OAI222 U516 ( .A(n1943), .B(n11037), .C(n1919), .D(n6594), .Q(n6961) );
  OAI222 U518 ( .A(n2279), .B(n11035), .C(n2255), .D(n6600), .Q(n6968) );
  OAI222 U519 ( .A(n2231), .B(n11033), .C(n2207), .D(n6602), .Q(n6967) );
  OAI222 U520 ( .A(n2183), .B(n11031), .C(n2159), .D(n6604), .Q(n6966) );
  OAI222 U521 ( .A(n2135), .B(n11029), .C(n2111), .D(n6606), .Q(n6965) );
  OAI222 U524 ( .A(n935), .B(n11027), .C(n911), .D(n6616), .Q(n6976) );
  OAI222 U525 ( .A(n887), .B(n11025), .C(n863), .D(n6618), .Q(n6975) );
  OAI222 U526 ( .A(n839), .B(n11023), .C(n815), .D(n6620), .Q(n6974) );
  OAI222 U527 ( .A(n791), .B(n11021), .C(n767), .D(n6622), .Q(n6973) );
  OAI222 U529 ( .A(n1127), .B(n11019), .C(n1103), .D(n6628), .Q(n6980) );
  OAI222 U530 ( .A(n1079), .B(n11017), .C(n1055), .D(n6630), .Q(n6979) );
  OAI222 U531 ( .A(n1031), .B(n11015), .C(n1007), .D(n6632), .Q(n6978) );
  OAI222 U532 ( .A(n983), .B(n11013), .C(n959), .D(n6634), .Q(n6977) );
  OAI222 U534 ( .A(n1319), .B(n11011), .C(n1295), .D(n6640), .Q(n6984) );
  OAI222 U535 ( .A(n1271), .B(n11009), .C(n1247), .D(n6642), .Q(n6983) );
  OAI222 U536 ( .A(n1223), .B(n11007), .C(n1199), .D(n6644), .Q(n6982) );
  OAI222 U537 ( .A(n1175), .B(n11005), .C(n1151), .D(n6646), .Q(n6981) );
  OAI222 U539 ( .A(n1511), .B(n11003), .C(n1487), .D(n6652), .Q(n6988) );
  OAI222 U540 ( .A(n1463), .B(n11001), .C(n1439), .D(n6654), .Q(n6987) );
  OAI222 U541 ( .A(n1415), .B(n10999), .C(n1391), .D(n6656), .Q(n6986) );
  OAI222 U542 ( .A(n1367), .B(n10997), .C(n1343), .D(n6658), .Q(n6985) );
  OAI222 U545 ( .A(n167), .B(n10995), .C(n143), .D(n6668), .Q(n6996) );
  OAI222 U546 ( .A(n119), .B(n10993), .C(n95), .D(n6670), .Q(n6995) );
  OAI222 U547 ( .A(n71), .B(n10991), .C(n47), .D(n6672), .Q(n6994) );
  OAI222 U548 ( .A(n23), .B(n10989), .C(n6143), .D(n6674), .Q(n6993) );
  OAI222 U550 ( .A(n359), .B(n10987), .C(n335), .D(n6680), .Q(n7000) );
  OAI222 U551 ( .A(n311), .B(n10985), .C(n287), .D(n6682), .Q(n6999) );
  OAI222 U552 ( .A(n263), .B(n10983), .C(n239), .D(n6684), .Q(n6998) );
  OAI222 U553 ( .A(n215), .B(n10981), .C(n191), .D(n6686), .Q(n6997) );
  OAI222 U555 ( .A(n551), .B(n10979), .C(n527), .D(n6692), .Q(n7004) );
  OAI222 U556 ( .A(n503), .B(n10977), .C(n479), .D(n6694), .Q(n7003) );
  OAI222 U557 ( .A(n455), .B(n10975), .C(n431), .D(n6696), .Q(n7002) );
  OAI222 U558 ( .A(n407), .B(n10973), .C(n383), .D(n6698), .Q(n7001) );
  OAI222 U560 ( .A(n743), .B(n10971), .C(n719), .D(n6704), .Q(n7008) );
  OAI222 U561 ( .A(n695), .B(n10969), .C(n671), .D(n6706), .Q(n7007) );
  OAI222 U562 ( .A(n647), .B(n10967), .C(n623), .D(n6708), .Q(n7006) );
  OAI222 U563 ( .A(n599), .B(n10965), .C(n575), .D(n6710), .Q(n7005) );
  OAI222 U567 ( .A(n5543), .B(n10963), .C(n5519), .D(n6724), .Q(n7020) );
  OAI222 U568 ( .A(n5495), .B(n10961), .C(n5471), .D(n6726), .Q(n7019) );
  OAI222 U569 ( .A(n5447), .B(n10959), .C(n5423), .D(n6728), .Q(n7018) );
  OAI222 U570 ( .A(n5399), .B(n10957), .C(n5375), .D(n6730), .Q(n7017) );
  OAI222 U572 ( .A(n5735), .B(n10955), .C(n5711), .D(n6736), .Q(n7024) );
  OAI222 U573 ( .A(n5687), .B(n10953), .C(n5663), .D(n6738), .Q(n7023) );
  OAI222 U574 ( .A(n5639), .B(n10951), .C(n5615), .D(n6740), .Q(n7022) );
  OAI222 U575 ( .A(n5591), .B(n10949), .C(n5567), .D(n6742), .Q(n7021) );
  OAI222 U577 ( .A(n5927), .B(n10947), .C(n5903), .D(n6748), .Q(n7028) );
  OAI222 U578 ( .A(n5879), .B(n10945), .C(n5855), .D(n6750), .Q(n7027) );
  OAI222 U579 ( .A(n5831), .B(n10943), .C(n5807), .D(n6752), .Q(n7026) );
  OAI222 U580 ( .A(n5783), .B(n10941), .C(n5759), .D(n6754), .Q(n7025) );
  OAI222 U582 ( .A(n6119), .B(n10939), .C(n6095), .D(n6760), .Q(n7032) );
  OAI222 U583 ( .A(n6071), .B(n10937), .C(n6047), .D(n6762), .Q(n7031) );
  OAI222 U584 ( .A(n6023), .B(n10935), .C(n5999), .D(n6764), .Q(n7030) );
  OAI222 U585 ( .A(n5975), .B(n10933), .C(n5951), .D(n6766), .Q(n7029) );
  OAI222 U588 ( .A(n4775), .B(n10931), .C(n4751), .D(n6776), .Q(n7040) );
  OAI222 U589 ( .A(n4727), .B(n10929), .C(n4703), .D(n6778), .Q(n7039) );
  OAI222 U590 ( .A(n4679), .B(n10927), .C(n4655), .D(n6780), .Q(n7038) );
  OAI222 U591 ( .A(n4631), .B(n10925), .C(n4607), .D(n6782), .Q(n7037) );
  OAI222 U593 ( .A(n4967), .B(n10923), .C(n4943), .D(n6788), .Q(n7044) );
  OAI222 U594 ( .A(n4919), .B(n10921), .C(n4895), .D(n6790), .Q(n7043) );
  OAI222 U595 ( .A(n4871), .B(n10919), .C(n4847), .D(n6792), .Q(n7042) );
  OAI222 U596 ( .A(n4823), .B(n10917), .C(n4799), .D(n6794), .Q(n7041) );
  OAI222 U598 ( .A(n5159), .B(n10915), .C(n5135), .D(n6800), .Q(n7048) );
  OAI222 U599 ( .A(n5111), .B(n10913), .C(n5087), .D(n6802), .Q(n7047) );
  OAI222 U600 ( .A(n5063), .B(n10911), .C(n5039), .D(n6804), .Q(n7046) );
  OAI222 U601 ( .A(n5015), .B(n10909), .C(n4991), .D(n6806), .Q(n7045) );
  OAI222 U603 ( .A(n5351), .B(n10907), .C(n5327), .D(n6812), .Q(n7052) );
  OAI222 U604 ( .A(n5303), .B(n10905), .C(n5279), .D(n6814), .Q(n7051) );
  OAI222 U605 ( .A(n5255), .B(n10903), .C(n5231), .D(n6816), .Q(n7050) );
  OAI222 U606 ( .A(n5207), .B(n10901), .C(n5183), .D(n6818), .Q(n7049) );
  OAI222 U609 ( .A(n4007), .B(n10899), .C(n3983), .D(n6828), .Q(n7060) );
  OAI222 U610 ( .A(n3959), .B(n10897), .C(n3935), .D(n6830), .Q(n7059) );
  OAI222 U611 ( .A(n3911), .B(n10895), .C(n3887), .D(n6832), .Q(n7058) );
  OAI222 U612 ( .A(n3863), .B(n10893), .C(n3839), .D(n6834), .Q(n7057) );
  OAI222 U614 ( .A(n4199), .B(n10891), .C(n4175), .D(n6840), .Q(n7064) );
  OAI222 U615 ( .A(n4151), .B(n10889), .C(n4127), .D(n6842), .Q(n7063) );
  OAI222 U616 ( .A(n4103), .B(n10887), .C(n4079), .D(n6844), .Q(n7062) );
  OAI222 U617 ( .A(n4055), .B(n10885), .C(n4031), .D(n6846), .Q(n7061) );
  OAI222 U619 ( .A(n4391), .B(n10883), .C(n4367), .D(n6852), .Q(n7068) );
  OAI222 U620 ( .A(n4343), .B(n10881), .C(n4319), .D(n6854), .Q(n7067) );
  OAI222 U621 ( .A(n4295), .B(n6191), .C(n4271), .D(n6856), .Q(n7066) );
  OAI222 U622 ( .A(n4247), .B(n6189), .C(n4223), .D(n6858), .Q(n7065) );
  OAI222 U624 ( .A(n4583), .B(n6187), .C(n4559), .D(n6864), .Q(n7072) );
  OAI222 U625 ( .A(n4535), .B(n6185), .C(n4511), .D(n6866), .Q(n7071) );
  OAI222 U626 ( .A(n4487), .B(n6183), .C(n4463), .D(n6868), .Q(n7070) );
  OAI222 U627 ( .A(n4439), .B(n6181), .C(n4415), .D(n6870), .Q(n7069) );
  OAI222 U630 ( .A(n3239), .B(n6179), .C(n3215), .D(n6880), .Q(n7080) );
  OAI222 U631 ( .A(n3191), .B(n6177), .C(n3167), .D(n6882), .Q(n7079) );
  OAI222 U632 ( .A(n3143), .B(n6175), .C(n3119), .D(n6884), .Q(n7078) );
  OAI222 U633 ( .A(n3095), .B(n6173), .C(n3071), .D(n6886), .Q(n7077) );
  OAI222 U635 ( .A(n3431), .B(n6171), .C(n3407), .D(n6892), .Q(n7084) );
  OAI222 U636 ( .A(n3383), .B(n6169), .C(n3359), .D(n6894), .Q(n7083) );
  OAI222 U637 ( .A(n3335), .B(n6167), .C(n3311), .D(n6896), .Q(n7082) );
  OAI222 U638 ( .A(n3287), .B(n6165), .C(n3263), .D(n6898), .Q(n7081) );
  OAI222 U640 ( .A(n3623), .B(n6163), .C(n3599), .D(n6904), .Q(n7088) );
  OAI222 U641 ( .A(n3575), .B(n6161), .C(n3551), .D(n6906), .Q(n7087) );
  OAI222 U642 ( .A(n3527), .B(n6159), .C(n3503), .D(n6908), .Q(n7086) );
  OAI222 U643 ( .A(n3479), .B(n6157), .C(n3455), .D(n6910), .Q(n7085) );
  OAI222 U645 ( .A(n3815), .B(n6155), .C(n3791), .D(n6916), .Q(n7092) );
  OAI222 U646 ( .A(n3767), .B(n6153), .C(n3743), .D(n6918), .Q(n7091) );
  OAI222 U647 ( .A(n3719), .B(n6151), .C(n3695), .D(n6920), .Q(n7090) );
  OAI222 U648 ( .A(n3671), .B(n6149), .C(n3647), .D(n6922), .Q(n7089) );
  OAI222 U653 ( .A(n2470), .B(n11091), .C(n2446), .D(n6512), .Q(n7106) );
  OAI222 U654 ( .A(n2422), .B(n11089), .C(n2398), .D(n6514), .Q(n7105) );
  OAI222 U655 ( .A(n2374), .B(n11087), .C(n2350), .D(n6516), .Q(n7104) );
  OAI222 U656 ( .A(n2326), .B(n11085), .C(n2302), .D(n6518), .Q(n7103) );
  OAI222 U658 ( .A(n2662), .B(n11083), .C(n2638), .D(n6524), .Q(n7110) );
  OAI222 U659 ( .A(n2614), .B(n11081), .C(n2590), .D(n6526), .Q(n7109) );
  OAI222 U660 ( .A(n2566), .B(n11079), .C(n2542), .D(n6528), .Q(n7108) );
  OAI222 U661 ( .A(n2518), .B(n11077), .C(n2494), .D(n6530), .Q(n7107) );
  OAI222 U663 ( .A(n2854), .B(n11075), .C(n2830), .D(n6536), .Q(n7114) );
  OAI222 U664 ( .A(n2806), .B(n11073), .C(n2782), .D(n6538), .Q(n7113) );
  OAI222 U665 ( .A(n2758), .B(n11071), .C(n2734), .D(n6540), .Q(n7112) );
  OAI222 U666 ( .A(n2710), .B(n11069), .C(n2686), .D(n6542), .Q(n7111) );
  OAI222 U668 ( .A(n3046), .B(n11067), .C(n3022), .D(n6548), .Q(n7118) );
  OAI222 U669 ( .A(n2998), .B(n11065), .C(n2974), .D(n6550), .Q(n7117) );
  OAI222 U670 ( .A(n2950), .B(n11063), .C(n2926), .D(n6552), .Q(n7116) );
  OAI222 U671 ( .A(n2902), .B(n11061), .C(n2878), .D(n6554), .Q(n7115) );
  OAI222 U674 ( .A(n1702), .B(n11059), .C(n1678), .D(n6564), .Q(n7126) );
  OAI222 U675 ( .A(n1654), .B(n11057), .C(n1630), .D(n6566), .Q(n7125) );
  OAI222 U676 ( .A(n1606), .B(n11055), .C(n1582), .D(n6568), .Q(n7124) );
  OAI222 U677 ( .A(n1558), .B(n11053), .C(n1534), .D(n6570), .Q(n7123) );
  OAI222 U679 ( .A(n1894), .B(n11051), .C(n1870), .D(n6576), .Q(n7130) );
  OAI222 U680 ( .A(n1846), .B(n11049), .C(n1822), .D(n6578), .Q(n7129) );
  OAI222 U681 ( .A(n1798), .B(n11047), .C(n1774), .D(n6580), .Q(n7128) );
  OAI222 U682 ( .A(n1750), .B(n11045), .C(n1726), .D(n6582), .Q(n7127) );
  OAI222 U684 ( .A(n2086), .B(n11043), .C(n2062), .D(n6588), .Q(n7134) );
  OAI222 U685 ( .A(n2038), .B(n11041), .C(n2014), .D(n6590), .Q(n7133) );
  OAI222 U686 ( .A(n1990), .B(n11039), .C(n1966), .D(n6592), .Q(n7132) );
  OAI222 U687 ( .A(n1942), .B(n11037), .C(n1918), .D(n6594), .Q(n7131) );
  OAI222 U689 ( .A(n2278), .B(n11035), .C(n2254), .D(n6600), .Q(n7138) );
  OAI222 U690 ( .A(n2230), .B(n11033), .C(n2206), .D(n6602), .Q(n7137) );
  OAI222 U691 ( .A(n2182), .B(n11031), .C(n2158), .D(n6604), .Q(n7136) );
  OAI222 U692 ( .A(n2134), .B(n11029), .C(n2110), .D(n6606), .Q(n7135) );
  OAI222 U695 ( .A(n934), .B(n11027), .C(n910), .D(n6616), .Q(n7146) );
  OAI222 U696 ( .A(n886), .B(n11025), .C(n862), .D(n6618), .Q(n7145) );
  OAI222 U697 ( .A(n838), .B(n11023), .C(n814), .D(n6620), .Q(n7144) );
  OAI222 U698 ( .A(n790), .B(n11021), .C(n766), .D(n6622), .Q(n7143) );
  OAI222 U700 ( .A(n1126), .B(n11019), .C(n1102), .D(n6628), .Q(n7150) );
  OAI222 U701 ( .A(n1078), .B(n11017), .C(n1054), .D(n6630), .Q(n7149) );
  OAI222 U702 ( .A(n1030), .B(n11015), .C(n1006), .D(n6632), .Q(n7148) );
  OAI222 U703 ( .A(n982), .B(n11013), .C(n958), .D(n6634), .Q(n7147) );
  OAI222 U705 ( .A(n1318), .B(n11011), .C(n1294), .D(n6640), .Q(n7154) );
  OAI222 U706 ( .A(n1270), .B(n11009), .C(n1246), .D(n6642), .Q(n7153) );
  OAI222 U707 ( .A(n1222), .B(n11007), .C(n1198), .D(n6644), .Q(n7152) );
  OAI222 U708 ( .A(n1174), .B(n11005), .C(n1150), .D(n6646), .Q(n7151) );
  OAI222 U710 ( .A(n1510), .B(n11003), .C(n1486), .D(n6652), .Q(n7158) );
  OAI222 U711 ( .A(n1462), .B(n11001), .C(n1438), .D(n6654), .Q(n7157) );
  OAI222 U712 ( .A(n1414), .B(n10999), .C(n1390), .D(n6656), .Q(n7156) );
  OAI222 U713 ( .A(n1366), .B(n10997), .C(n1342), .D(n6658), .Q(n7155) );
  OAI222 U716 ( .A(n166), .B(n10995), .C(n142), .D(n6668), .Q(n7166) );
  OAI222 U717 ( .A(n118), .B(n10993), .C(n94), .D(n6670), .Q(n7165) );
  OAI222 U718 ( .A(n70), .B(n10991), .C(n46), .D(n6672), .Q(n7164) );
  OAI222 U719 ( .A(n22), .B(n10989), .C(n6142), .D(n6674), .Q(n7163) );
  OAI222 U721 ( .A(n358), .B(n10987), .C(n334), .D(n6680), .Q(n7170) );
  OAI222 U722 ( .A(n310), .B(n10985), .C(n286), .D(n6682), .Q(n7169) );
  OAI222 U723 ( .A(n262), .B(n10983), .C(n238), .D(n6684), .Q(n7168) );
  OAI222 U724 ( .A(n214), .B(n10981), .C(n190), .D(n6686), .Q(n7167) );
  OAI222 U726 ( .A(n550), .B(n10979), .C(n526), .D(n6692), .Q(n7174) );
  OAI222 U727 ( .A(n502), .B(n10977), .C(n478), .D(n6694), .Q(n7173) );
  OAI222 U728 ( .A(n454), .B(n10975), .C(n430), .D(n6696), .Q(n7172) );
  OAI222 U729 ( .A(n406), .B(n10973), .C(n382), .D(n6698), .Q(n7171) );
  OAI222 U731 ( .A(n742), .B(n10971), .C(n718), .D(n6704), .Q(n7178) );
  OAI222 U732 ( .A(n694), .B(n10969), .C(n670), .D(n6706), .Q(n7177) );
  OAI222 U733 ( .A(n646), .B(n10967), .C(n622), .D(n6708), .Q(n7176) );
  OAI222 U734 ( .A(n598), .B(n10965), .C(n574), .D(n6710), .Q(n7175) );
  OAI222 U738 ( .A(n5542), .B(n10963), .C(n5518), .D(n6724), .Q(n7190) );
  OAI222 U739 ( .A(n5494), .B(n10961), .C(n5470), .D(n6726), .Q(n7189) );
  OAI222 U740 ( .A(n5446), .B(n10959), .C(n5422), .D(n6728), .Q(n7188) );
  OAI222 U741 ( .A(n5398), .B(n10957), .C(n5374), .D(n6730), .Q(n7187) );
  OAI222 U743 ( .A(n5734), .B(n10955), .C(n5710), .D(n6736), .Q(n7194) );
  OAI222 U744 ( .A(n5686), .B(n10953), .C(n5662), .D(n6738), .Q(n7193) );
  OAI222 U745 ( .A(n5638), .B(n10951), .C(n5614), .D(n6740), .Q(n7192) );
  OAI222 U746 ( .A(n5590), .B(n10949), .C(n5566), .D(n6742), .Q(n7191) );
  OAI222 U748 ( .A(n5926), .B(n10947), .C(n5902), .D(n6748), .Q(n7198) );
  OAI222 U749 ( .A(n5878), .B(n10945), .C(n5854), .D(n6750), .Q(n7197) );
  OAI222 U750 ( .A(n5830), .B(n10943), .C(n5806), .D(n6752), .Q(n7196) );
  OAI222 U751 ( .A(n5782), .B(n10941), .C(n5758), .D(n6754), .Q(n7195) );
  OAI222 U753 ( .A(n6118), .B(n10939), .C(n6094), .D(n6760), .Q(n7202) );
  OAI222 U754 ( .A(n6070), .B(n10937), .C(n6046), .D(n6762), .Q(n7201) );
  OAI222 U755 ( .A(n6022), .B(n10935), .C(n5998), .D(n6764), .Q(n7200) );
  OAI222 U756 ( .A(n5974), .B(n10933), .C(n5950), .D(n6766), .Q(n7199) );
  OAI222 U759 ( .A(n4774), .B(n10931), .C(n4750), .D(n6776), .Q(n7210) );
  OAI222 U760 ( .A(n4726), .B(n10929), .C(n4702), .D(n6778), .Q(n7209) );
  OAI222 U761 ( .A(n4678), .B(n10927), .C(n4654), .D(n6780), .Q(n7208) );
  OAI222 U762 ( .A(n4630), .B(n10925), .C(n4606), .D(n6782), .Q(n7207) );
  OAI222 U764 ( .A(n4966), .B(n10923), .C(n4942), .D(n6788), .Q(n7214) );
  OAI222 U765 ( .A(n4918), .B(n10921), .C(n4894), .D(n6790), .Q(n7213) );
  OAI222 U766 ( .A(n4870), .B(n10919), .C(n4846), .D(n6792), .Q(n7212) );
  OAI222 U767 ( .A(n4822), .B(n10917), .C(n4798), .D(n6794), .Q(n7211) );
  OAI222 U769 ( .A(n5158), .B(n10915), .C(n5134), .D(n6800), .Q(n7218) );
  OAI222 U770 ( .A(n5110), .B(n10913), .C(n5086), .D(n6802), .Q(n7217) );
  OAI222 U771 ( .A(n5062), .B(n10911), .C(n5038), .D(n6804), .Q(n7216) );
  OAI222 U772 ( .A(n5014), .B(n10909), .C(n4990), .D(n6806), .Q(n7215) );
  OAI222 U774 ( .A(n5350), .B(n10907), .C(n5326), .D(n6812), .Q(n7222) );
  OAI222 U775 ( .A(n5302), .B(n10905), .C(n5278), .D(n6814), .Q(n7221) );
  OAI222 U776 ( .A(n5254), .B(n10903), .C(n5230), .D(n6816), .Q(n7220) );
  OAI222 U777 ( .A(n5206), .B(n10901), .C(n5182), .D(n6818), .Q(n7219) );
  OAI222 U780 ( .A(n4006), .B(n10899), .C(n3982), .D(n6828), .Q(n7230) );
  OAI222 U781 ( .A(n3958), .B(n10897), .C(n3934), .D(n6830), .Q(n7229) );
  OAI222 U782 ( .A(n3910), .B(n10895), .C(n3886), .D(n6832), .Q(n7228) );
  OAI222 U783 ( .A(n3862), .B(n10893), .C(n3838), .D(n6834), .Q(n7227) );
  OAI222 U785 ( .A(n4198), .B(n10891), .C(n4174), .D(n6840), .Q(n7234) );
  OAI222 U786 ( .A(n4150), .B(n10889), .C(n4126), .D(n6842), .Q(n7233) );
  OAI222 U787 ( .A(n4102), .B(n10887), .C(n4078), .D(n6844), .Q(n7232) );
  OAI222 U788 ( .A(n4054), .B(n10885), .C(n4030), .D(n6846), .Q(n7231) );
  OAI222 U790 ( .A(n4390), .B(n10883), .C(n4366), .D(n6852), .Q(n7238) );
  OAI222 U791 ( .A(n4342), .B(n10881), .C(n4318), .D(n6854), .Q(n7237) );
  OAI222 U792 ( .A(n4294), .B(n6191), .C(n4270), .D(n6856), .Q(n7236) );
  OAI222 U793 ( .A(n4246), .B(n6189), .C(n4222), .D(n6858), .Q(n7235) );
  OAI222 U795 ( .A(n4582), .B(n6187), .C(n4558), .D(n6864), .Q(n7242) );
  OAI222 U796 ( .A(n4534), .B(n6185), .C(n4510), .D(n6866), .Q(n7241) );
  OAI222 U797 ( .A(n4486), .B(n6183), .C(n4462), .D(n6868), .Q(n7240) );
  OAI222 U798 ( .A(n4438), .B(n6181), .C(n4414), .D(n6870), .Q(n7239) );
  OAI222 U801 ( .A(n3238), .B(n6179), .C(n3214), .D(n6880), .Q(n7250) );
  OAI222 U802 ( .A(n3190), .B(n6177), .C(n3166), .D(n6882), .Q(n7249) );
  OAI222 U803 ( .A(n3142), .B(n6175), .C(n3118), .D(n6884), .Q(n7248) );
  OAI222 U804 ( .A(n3094), .B(n6173), .C(n3070), .D(n6886), .Q(n7247) );
  OAI222 U806 ( .A(n3430), .B(n6171), .C(n3406), .D(n6892), .Q(n7254) );
  OAI222 U807 ( .A(n3382), .B(n6169), .C(n3358), .D(n6894), .Q(n7253) );
  OAI222 U808 ( .A(n3334), .B(n6167), .C(n3310), .D(n6896), .Q(n7252) );
  OAI222 U809 ( .A(n3286), .B(n6165), .C(n3262), .D(n6898), .Q(n7251) );
  OAI222 U811 ( .A(n3622), .B(n6163), .C(n3598), .D(n6904), .Q(n7258) );
  OAI222 U812 ( .A(n3574), .B(n6161), .C(n3550), .D(n6906), .Q(n7257) );
  OAI222 U813 ( .A(n3526), .B(n6159), .C(n3502), .D(n6908), .Q(n7256) );
  OAI222 U814 ( .A(n3478), .B(n6157), .C(n3454), .D(n6910), .Q(n7255) );
  OAI222 U816 ( .A(n3814), .B(n6155), .C(n3790), .D(n6916), .Q(n7262) );
  OAI222 U817 ( .A(n3766), .B(n6153), .C(n3742), .D(n6918), .Q(n7261) );
  OAI222 U818 ( .A(n3718), .B(n6151), .C(n3694), .D(n6920), .Q(n7260) );
  OAI222 U819 ( .A(n3670), .B(n6149), .C(n3646), .D(n6922), .Q(n7259) );
  OAI222 U824 ( .A(n2469), .B(n11091), .C(n2445), .D(n6512), .Q(n7276) );
  OAI222 U825 ( .A(n2421), .B(n11089), .C(n2397), .D(n6514), .Q(n7275) );
  OAI222 U826 ( .A(n2373), .B(n11087), .C(n2349), .D(n6516), .Q(n7274) );
  OAI222 U827 ( .A(n2325), .B(n11085), .C(n2301), .D(n6518), .Q(n7273) );
  OAI222 U829 ( .A(n2661), .B(n11083), .C(n2637), .D(n6524), .Q(n7280) );
  OAI222 U830 ( .A(n2613), .B(n11081), .C(n2589), .D(n6526), .Q(n7279) );
  OAI222 U831 ( .A(n2565), .B(n11079), .C(n2541), .D(n6528), .Q(n7278) );
  OAI222 U832 ( .A(n2517), .B(n11077), .C(n2493), .D(n6530), .Q(n7277) );
  OAI222 U834 ( .A(n2853), .B(n11075), .C(n2829), .D(n6536), .Q(n7284) );
  OAI222 U835 ( .A(n2805), .B(n11073), .C(n2781), .D(n6538), .Q(n7283) );
  OAI222 U836 ( .A(n2757), .B(n11071), .C(n2733), .D(n6540), .Q(n7282) );
  OAI222 U837 ( .A(n2709), .B(n11069), .C(n2685), .D(n6542), .Q(n7281) );
  OAI222 U839 ( .A(n3045), .B(n11067), .C(n3021), .D(n6548), .Q(n7288) );
  OAI222 U840 ( .A(n2997), .B(n11065), .C(n2973), .D(n6550), .Q(n7287) );
  OAI222 U841 ( .A(n2949), .B(n11063), .C(n2925), .D(n6552), .Q(n7286) );
  OAI222 U842 ( .A(n2901), .B(n11061), .C(n2877), .D(n6554), .Q(n7285) );
  OAI222 U845 ( .A(n1701), .B(n11059), .C(n1677), .D(n6564), .Q(n7296) );
  OAI222 U846 ( .A(n1653), .B(n11057), .C(n1629), .D(n6566), .Q(n7295) );
  OAI222 U847 ( .A(n1605), .B(n11055), .C(n1581), .D(n6568), .Q(n7294) );
  OAI222 U848 ( .A(n1557), .B(n11053), .C(n1533), .D(n6570), .Q(n7293) );
  OAI222 U850 ( .A(n1893), .B(n11051), .C(n1869), .D(n6576), .Q(n7300) );
  OAI222 U851 ( .A(n1845), .B(n11049), .C(n1821), .D(n6578), .Q(n7299) );
  OAI222 U852 ( .A(n1797), .B(n11047), .C(n1773), .D(n6580), .Q(n7298) );
  OAI222 U853 ( .A(n1749), .B(n11045), .C(n1725), .D(n6582), .Q(n7297) );
  OAI222 U855 ( .A(n2085), .B(n11043), .C(n2061), .D(n6588), .Q(n7304) );
  OAI222 U856 ( .A(n2037), .B(n11041), .C(n2013), .D(n6590), .Q(n7303) );
  OAI222 U857 ( .A(n1989), .B(n11039), .C(n1965), .D(n6592), .Q(n7302) );
  OAI222 U858 ( .A(n1941), .B(n11037), .C(n1917), .D(n6594), .Q(n7301) );
  OAI222 U860 ( .A(n2277), .B(n11035), .C(n2253), .D(n6600), .Q(n7308) );
  OAI222 U861 ( .A(n2229), .B(n11033), .C(n2205), .D(n6602), .Q(n7307) );
  OAI222 U862 ( .A(n2181), .B(n11031), .C(n2157), .D(n6604), .Q(n7306) );
  OAI222 U863 ( .A(n2133), .B(n11029), .C(n2109), .D(n6606), .Q(n7305) );
  OAI222 U866 ( .A(n933), .B(n11027), .C(n909), .D(n6616), .Q(n7316) );
  OAI222 U867 ( .A(n885), .B(n11025), .C(n861), .D(n6618), .Q(n7315) );
  OAI222 U868 ( .A(n837), .B(n11023), .C(n813), .D(n6620), .Q(n7314) );
  OAI222 U869 ( .A(n789), .B(n11021), .C(n765), .D(n6622), .Q(n7313) );
  OAI222 U871 ( .A(n1125), .B(n11019), .C(n1101), .D(n6628), .Q(n7320) );
  OAI222 U872 ( .A(n1077), .B(n11017), .C(n1053), .D(n6630), .Q(n7319) );
  OAI222 U873 ( .A(n1029), .B(n11015), .C(n1005), .D(n6632), .Q(n7318) );
  OAI222 U874 ( .A(n981), .B(n11013), .C(n957), .D(n6634), .Q(n7317) );
  OAI222 U876 ( .A(n1317), .B(n11011), .C(n1293), .D(n6640), .Q(n7324) );
  OAI222 U877 ( .A(n1269), .B(n11009), .C(n1245), .D(n6642), .Q(n7323) );
  OAI222 U878 ( .A(n1221), .B(n11007), .C(n1197), .D(n6644), .Q(n7322) );
  OAI222 U879 ( .A(n1173), .B(n11005), .C(n1149), .D(n6646), .Q(n7321) );
  OAI222 U881 ( .A(n1509), .B(n11003), .C(n1485), .D(n6652), .Q(n7328) );
  OAI222 U882 ( .A(n1461), .B(n11001), .C(n1437), .D(n6654), .Q(n7327) );
  OAI222 U883 ( .A(n1413), .B(n10999), .C(n1389), .D(n6656), .Q(n7326) );
  OAI222 U884 ( .A(n1365), .B(n10997), .C(n1341), .D(n6658), .Q(n7325) );
  OAI222 U887 ( .A(n165), .B(n10995), .C(n141), .D(n6668), .Q(n7336) );
  OAI222 U888 ( .A(n117), .B(n10993), .C(n93), .D(n6670), .Q(n7335) );
  OAI222 U889 ( .A(n69), .B(n10991), .C(n45), .D(n6672), .Q(n7334) );
  OAI222 U890 ( .A(n21), .B(n10989), .C(n6141), .D(n6674), .Q(n7333) );
  OAI222 U892 ( .A(n357), .B(n10987), .C(n333), .D(n6680), .Q(n7340) );
  OAI222 U893 ( .A(n309), .B(n10985), .C(n285), .D(n6682), .Q(n7339) );
  OAI222 U894 ( .A(n261), .B(n10983), .C(n237), .D(n6684), .Q(n7338) );
  OAI222 U895 ( .A(n213), .B(n10981), .C(n189), .D(n6686), .Q(n7337) );
  OAI222 U897 ( .A(n549), .B(n10979), .C(n525), .D(n6692), .Q(n7344) );
  OAI222 U898 ( .A(n501), .B(n10977), .C(n477), .D(n6694), .Q(n7343) );
  OAI222 U899 ( .A(n453), .B(n10975), .C(n429), .D(n6696), .Q(n7342) );
  OAI222 U900 ( .A(n405), .B(n10973), .C(n381), .D(n6698), .Q(n7341) );
  OAI222 U902 ( .A(n741), .B(n10971), .C(n717), .D(n6704), .Q(n7348) );
  OAI222 U903 ( .A(n693), .B(n10969), .C(n669), .D(n6706), .Q(n7347) );
  OAI222 U904 ( .A(n645), .B(n10967), .C(n621), .D(n6708), .Q(n7346) );
  OAI222 U905 ( .A(n597), .B(n10965), .C(n573), .D(n6710), .Q(n7345) );
  OAI222 U909 ( .A(n5541), .B(n10963), .C(n5517), .D(n6724), .Q(n7360) );
  OAI222 U910 ( .A(n5493), .B(n10961), .C(n5469), .D(n6726), .Q(n7359) );
  OAI222 U911 ( .A(n5445), .B(n10959), .C(n5421), .D(n6728), .Q(n7358) );
  OAI222 U912 ( .A(n5397), .B(n10957), .C(n5373), .D(n6730), .Q(n7357) );
  OAI222 U914 ( .A(n5733), .B(n10955), .C(n5709), .D(n6736), .Q(n7364) );
  OAI222 U915 ( .A(n5685), .B(n10953), .C(n5661), .D(n6738), .Q(n7363) );
  OAI222 U916 ( .A(n5637), .B(n10951), .C(n5613), .D(n6740), .Q(n7362) );
  OAI222 U917 ( .A(n5589), .B(n10949), .C(n5565), .D(n6742), .Q(n7361) );
  OAI222 U919 ( .A(n5925), .B(n10947), .C(n5901), .D(n6748), .Q(n7368) );
  OAI222 U920 ( .A(n5877), .B(n10945), .C(n5853), .D(n6750), .Q(n7367) );
  OAI222 U921 ( .A(n5829), .B(n10943), .C(n5805), .D(n6752), .Q(n7366) );
  OAI222 U922 ( .A(n5781), .B(n10941), .C(n5757), .D(n6754), .Q(n7365) );
  OAI222 U924 ( .A(n6117), .B(n10939), .C(n6093), .D(n6760), .Q(n7372) );
  OAI222 U925 ( .A(n6069), .B(n10937), .C(n6045), .D(n6762), .Q(n7371) );
  OAI222 U926 ( .A(n6021), .B(n10935), .C(n5997), .D(n6764), .Q(n7370) );
  OAI222 U927 ( .A(n5973), .B(n10933), .C(n5949), .D(n6766), .Q(n7369) );
  OAI222 U930 ( .A(n4773), .B(n10931), .C(n4749), .D(n6776), .Q(n7380) );
  OAI222 U931 ( .A(n4725), .B(n10929), .C(n4701), .D(n6778), .Q(n7379) );
  OAI222 U932 ( .A(n4677), .B(n10927), .C(n4653), .D(n6780), .Q(n7378) );
  OAI222 U933 ( .A(n4629), .B(n10925), .C(n4605), .D(n6782), .Q(n7377) );
  OAI222 U935 ( .A(n4965), .B(n10923), .C(n4941), .D(n6788), .Q(n7384) );
  OAI222 U936 ( .A(n4917), .B(n10921), .C(n4893), .D(n6790), .Q(n7383) );
  OAI222 U937 ( .A(n4869), .B(n10919), .C(n4845), .D(n6792), .Q(n7382) );
  OAI222 U938 ( .A(n4821), .B(n10917), .C(n4797), .D(n6794), .Q(n7381) );
  OAI222 U940 ( .A(n5157), .B(n10915), .C(n5133), .D(n6800), .Q(n7388) );
  OAI222 U941 ( .A(n5109), .B(n10913), .C(n5085), .D(n6802), .Q(n7387) );
  OAI222 U942 ( .A(n5061), .B(n10911), .C(n5037), .D(n6804), .Q(n7386) );
  OAI222 U943 ( .A(n5013), .B(n10909), .C(n4989), .D(n6806), .Q(n7385) );
  OAI222 U945 ( .A(n5349), .B(n10907), .C(n5325), .D(n6812), .Q(n7392) );
  OAI222 U946 ( .A(n5301), .B(n10905), .C(n5277), .D(n6814), .Q(n7391) );
  OAI222 U947 ( .A(n5253), .B(n10903), .C(n5229), .D(n6816), .Q(n7390) );
  OAI222 U948 ( .A(n5205), .B(n10901), .C(n5181), .D(n6818), .Q(n7389) );
  OAI222 U951 ( .A(n4005), .B(n10899), .C(n3981), .D(n6828), .Q(n7400) );
  OAI222 U952 ( .A(n3957), .B(n10897), .C(n3933), .D(n6830), .Q(n7399) );
  OAI222 U953 ( .A(n3909), .B(n10895), .C(n3885), .D(n6832), .Q(n7398) );
  OAI222 U954 ( .A(n3861), .B(n10893), .C(n3837), .D(n6834), .Q(n7397) );
  OAI222 U956 ( .A(n4197), .B(n10891), .C(n4173), .D(n6840), .Q(n7404) );
  OAI222 U957 ( .A(n4149), .B(n10889), .C(n4125), .D(n6842), .Q(n7403) );
  OAI222 U958 ( .A(n4101), .B(n10887), .C(n4077), .D(n6844), .Q(n7402) );
  OAI222 U959 ( .A(n4053), .B(n10885), .C(n4029), .D(n6846), .Q(n7401) );
  OAI222 U961 ( .A(n4389), .B(n10883), .C(n4365), .D(n6852), .Q(n7408) );
  OAI222 U962 ( .A(n4341), .B(n10881), .C(n4317), .D(n6854), .Q(n7407) );
  OAI222 U963 ( .A(n4293), .B(n6191), .C(n4269), .D(n6856), .Q(n7406) );
  OAI222 U964 ( .A(n4245), .B(n6189), .C(n4221), .D(n6858), .Q(n7405) );
  OAI222 U966 ( .A(n4581), .B(n6187), .C(n4557), .D(n6864), .Q(n7412) );
  OAI222 U967 ( .A(n4533), .B(n6185), .C(n4509), .D(n6866), .Q(n7411) );
  OAI222 U968 ( .A(n4485), .B(n6183), .C(n4461), .D(n6868), .Q(n7410) );
  OAI222 U969 ( .A(n4437), .B(n6181), .C(n4413), .D(n6870), .Q(n7409) );
  OAI222 U972 ( .A(n3237), .B(n6179), .C(n3213), .D(n6880), .Q(n7420) );
  OAI222 U973 ( .A(n3189), .B(n6177), .C(n3165), .D(n6882), .Q(n7419) );
  OAI222 U974 ( .A(n3141), .B(n6175), .C(n3117), .D(n6884), .Q(n7418) );
  OAI222 U975 ( .A(n3093), .B(n6173), .C(n3069), .D(n6886), .Q(n7417) );
  OAI222 U977 ( .A(n3429), .B(n6171), .C(n3405), .D(n6892), .Q(n7424) );
  OAI222 U978 ( .A(n3381), .B(n6169), .C(n3357), .D(n6894), .Q(n7423) );
  OAI222 U979 ( .A(n3333), .B(n6167), .C(n3309), .D(n6896), .Q(n7422) );
  OAI222 U980 ( .A(n3285), .B(n6165), .C(n3261), .D(n6898), .Q(n7421) );
  OAI222 U982 ( .A(n3621), .B(n6163), .C(n3597), .D(n6904), .Q(n7428) );
  OAI222 U983 ( .A(n3573), .B(n6161), .C(n3549), .D(n6906), .Q(n7427) );
  OAI222 U984 ( .A(n3525), .B(n6159), .C(n3501), .D(n6908), .Q(n7426) );
  OAI222 U985 ( .A(n3477), .B(n6157), .C(n3453), .D(n6910), .Q(n7425) );
  OAI222 U987 ( .A(n3813), .B(n6155), .C(n3789), .D(n6916), .Q(n7432) );
  OAI222 U988 ( .A(n3765), .B(n6153), .C(n3741), .D(n6918), .Q(n7431) );
  OAI222 U989 ( .A(n3717), .B(n6151), .C(n3693), .D(n6920), .Q(n7430) );
  OAI222 U990 ( .A(n3669), .B(n6149), .C(n3645), .D(n6922), .Q(n7429) );
  OAI222 U995 ( .A(n2468), .B(n11091), .C(n2444), .D(n6512), .Q(n7446) );
  OAI222 U996 ( .A(n2420), .B(n11089), .C(n2396), .D(n6514), .Q(n7445) );
  OAI222 U997 ( .A(n2372), .B(n11087), .C(n2348), .D(n6516), .Q(n7444) );
  OAI222 U998 ( .A(n2324), .B(n11085), .C(n2300), .D(n6518), .Q(n7443) );
  OAI222 U1000 ( .A(n2660), .B(n11083), .C(n2636), .D(n6524), .Q(n7450) );
  OAI222 U1001 ( .A(n2612), .B(n11081), .C(n2588), .D(n6526), .Q(n7449) );
  OAI222 U1002 ( .A(n2564), .B(n11079), .C(n2540), .D(n6528), .Q(n7448) );
  OAI222 U1003 ( .A(n2516), .B(n11077), .C(n2492), .D(n6530), .Q(n7447) );
  OAI222 U1005 ( .A(n2852), .B(n11075), .C(n2828), .D(n6536), .Q(n7454) );
  OAI222 U1006 ( .A(n2804), .B(n11073), .C(n2780), .D(n6538), .Q(n7453) );
  OAI222 U1007 ( .A(n2756), .B(n11071), .C(n2732), .D(n6540), .Q(n7452) );
  OAI222 U1008 ( .A(n2708), .B(n11069), .C(n2684), .D(n6542), .Q(n7451) );
  OAI222 U1010 ( .A(n3044), .B(n11067), .C(n3020), .D(n6548), .Q(n7458) );
  OAI222 U1011 ( .A(n2996), .B(n11065), .C(n2972), .D(n6550), .Q(n7457) );
  OAI222 U1012 ( .A(n2948), .B(n11063), .C(n2924), .D(n6552), .Q(n7456) );
  OAI222 U1013 ( .A(n2900), .B(n11061), .C(n2876), .D(n6554), .Q(n7455) );
  OAI222 U1016 ( .A(n1700), .B(n11059), .C(n1676), .D(n6564), .Q(n7466) );
  OAI222 U1017 ( .A(n1652), .B(n11057), .C(n1628), .D(n6566), .Q(n7465) );
  OAI222 U1018 ( .A(n1604), .B(n11055), .C(n1580), .D(n6568), .Q(n7464) );
  OAI222 U1019 ( .A(n1556), .B(n11053), .C(n1532), .D(n6570), .Q(n7463) );
  OAI222 U1021 ( .A(n1892), .B(n11051), .C(n1868), .D(n6576), .Q(n7470) );
  OAI222 U1022 ( .A(n1844), .B(n11049), .C(n1820), .D(n6578), .Q(n7469) );
  OAI222 U1023 ( .A(n1796), .B(n11047), .C(n1772), .D(n6580), .Q(n7468) );
  OAI222 U1024 ( .A(n1748), .B(n11045), .C(n1724), .D(n6582), .Q(n7467) );
  OAI222 U1026 ( .A(n2084), .B(n11043), .C(n2060), .D(n6588), .Q(n7474) );
  OAI222 U1027 ( .A(n2036), .B(n11041), .C(n2012), .D(n6590), .Q(n7473) );
  OAI222 U1028 ( .A(n1988), .B(n11039), .C(n1964), .D(n6592), .Q(n7472) );
  OAI222 U1029 ( .A(n1940), .B(n11037), .C(n1916), .D(n6594), .Q(n7471) );
  OAI222 U1031 ( .A(n2276), .B(n11035), .C(n2252), .D(n6600), .Q(n7478) );
  OAI222 U1032 ( .A(n2228), .B(n11033), .C(n2204), .D(n6602), .Q(n7477) );
  OAI222 U1033 ( .A(n2180), .B(n11031), .C(n2156), .D(n6604), .Q(n7476) );
  OAI222 U1034 ( .A(n2132), .B(n11029), .C(n2108), .D(n6606), .Q(n7475) );
  OAI222 U1037 ( .A(n932), .B(n11027), .C(n908), .D(n6616), .Q(n7486) );
  OAI222 U1038 ( .A(n884), .B(n11025), .C(n860), .D(n6618), .Q(n7485) );
  OAI222 U1039 ( .A(n836), .B(n11023), .C(n812), .D(n6620), .Q(n7484) );
  OAI222 U1040 ( .A(n788), .B(n11021), .C(n764), .D(n6622), .Q(n7483) );
  OAI222 U1042 ( .A(n1124), .B(n11019), .C(n1100), .D(n6628), .Q(n7490) );
  OAI222 U1043 ( .A(n1076), .B(n11017), .C(n1052), .D(n6630), .Q(n7489) );
  OAI222 U1044 ( .A(n1028), .B(n11015), .C(n1004), .D(n6632), .Q(n7488) );
  OAI222 U1045 ( .A(n980), .B(n11013), .C(n956), .D(n6634), .Q(n7487) );
  OAI222 U1047 ( .A(n1316), .B(n11011), .C(n1292), .D(n6640), .Q(n7494) );
  OAI222 U1048 ( .A(n1268), .B(n11009), .C(n1244), .D(n6642), .Q(n7493) );
  OAI222 U1049 ( .A(n1220), .B(n11007), .C(n1196), .D(n6644), .Q(n7492) );
  OAI222 U1050 ( .A(n1172), .B(n11005), .C(n1148), .D(n6646), .Q(n7491) );
  OAI222 U1052 ( .A(n1508), .B(n11003), .C(n1484), .D(n6652), .Q(n7498) );
  OAI222 U1053 ( .A(n1460), .B(n11001), .C(n1436), .D(n6654), .Q(n7497) );
  OAI222 U1054 ( .A(n1412), .B(n10999), .C(n1388), .D(n6656), .Q(n7496) );
  OAI222 U1055 ( .A(n1364), .B(n10997), .C(n1340), .D(n6658), .Q(n7495) );
  OAI222 U1058 ( .A(n164), .B(n10995), .C(n140), .D(n6668), .Q(n7506) );
  OAI222 U1059 ( .A(n116), .B(n10993), .C(n92), .D(n6670), .Q(n7505) );
  OAI222 U1060 ( .A(n68), .B(n10991), .C(n44), .D(n6672), .Q(n7504) );
  OAI222 U1061 ( .A(n20), .B(n10989), .C(n6140), .D(n6674), .Q(n7503) );
  OAI222 U1063 ( .A(n356), .B(n10987), .C(n332), .D(n6680), .Q(n7510) );
  OAI222 U1064 ( .A(n308), .B(n10985), .C(n284), .D(n6682), .Q(n7509) );
  OAI222 U1065 ( .A(n260), .B(n10983), .C(n236), .D(n6684), .Q(n7508) );
  OAI222 U1066 ( .A(n212), .B(n10981), .C(n188), .D(n6686), .Q(n7507) );
  OAI222 U1068 ( .A(n548), .B(n10979), .C(n524), .D(n6692), .Q(n7514) );
  OAI222 U1069 ( .A(n500), .B(n10977), .C(n476), .D(n6694), .Q(n7513) );
  OAI222 U1070 ( .A(n452), .B(n10975), .C(n428), .D(n6696), .Q(n7512) );
  OAI222 U1071 ( .A(n404), .B(n10973), .C(n380), .D(n6698), .Q(n7511) );
  OAI222 U1073 ( .A(n740), .B(n10971), .C(n716), .D(n6704), .Q(n7518) );
  OAI222 U1074 ( .A(n692), .B(n10969), .C(n668), .D(n6706), .Q(n7517) );
  OAI222 U1075 ( .A(n644), .B(n10967), .C(n620), .D(n6708), .Q(n7516) );
  OAI222 U1076 ( .A(n596), .B(n10965), .C(n572), .D(n6710), .Q(n7515) );
  OAI222 U1080 ( .A(n5540), .B(n10963), .C(n5516), .D(n6724), .Q(n7530) );
  OAI222 U1081 ( .A(n5492), .B(n10961), .C(n5468), .D(n6726), .Q(n7529) );
  OAI222 U1082 ( .A(n5444), .B(n10959), .C(n5420), .D(n6728), .Q(n7528) );
  OAI222 U1083 ( .A(n5396), .B(n10957), .C(n5372), .D(n6730), .Q(n7527) );
  OAI222 U1085 ( .A(n5732), .B(n10955), .C(n5708), .D(n6736), .Q(n7534) );
  OAI222 U1086 ( .A(n5684), .B(n10953), .C(n5660), .D(n6738), .Q(n7533) );
  OAI222 U1087 ( .A(n5636), .B(n10951), .C(n5612), .D(n6740), .Q(n7532) );
  OAI222 U1088 ( .A(n5588), .B(n10949), .C(n5564), .D(n6742), .Q(n7531) );
  OAI222 U1090 ( .A(n5924), .B(n10947), .C(n5900), .D(n6748), .Q(n7538) );
  OAI222 U1091 ( .A(n5876), .B(n10945), .C(n5852), .D(n6750), .Q(n7537) );
  OAI222 U1092 ( .A(n5828), .B(n10943), .C(n5804), .D(n6752), .Q(n7536) );
  OAI222 U1093 ( .A(n5780), .B(n10941), .C(n5756), .D(n6754), .Q(n7535) );
  OAI222 U1095 ( .A(n6116), .B(n10939), .C(n6092), .D(n6760), .Q(n7542) );
  OAI222 U1096 ( .A(n6068), .B(n10937), .C(n6044), .D(n6762), .Q(n7541) );
  OAI222 U1097 ( .A(n6020), .B(n10935), .C(n5996), .D(n6764), .Q(n7540) );
  OAI222 U1098 ( .A(n5972), .B(n10933), .C(n5948), .D(n6766), .Q(n7539) );
  OAI222 U1101 ( .A(n4772), .B(n10931), .C(n4748), .D(n6776), .Q(n7550) );
  OAI222 U1102 ( .A(n4724), .B(n10929), .C(n4700), .D(n6778), .Q(n7549) );
  OAI222 U1103 ( .A(n4676), .B(n10927), .C(n4652), .D(n6780), .Q(n7548) );
  OAI222 U1104 ( .A(n4628), .B(n10925), .C(n4604), .D(n6782), .Q(n7547) );
  OAI222 U1106 ( .A(n4964), .B(n10923), .C(n4940), .D(n6788), .Q(n7554) );
  OAI222 U1107 ( .A(n4916), .B(n10921), .C(n4892), .D(n6790), .Q(n7553) );
  OAI222 U1108 ( .A(n4868), .B(n10919), .C(n4844), .D(n6792), .Q(n7552) );
  OAI222 U1109 ( .A(n4820), .B(n10917), .C(n4796), .D(n6794), .Q(n7551) );
  OAI222 U1111 ( .A(n5156), .B(n10915), .C(n5132), .D(n6800), .Q(n7558) );
  OAI222 U1112 ( .A(n5108), .B(n10913), .C(n5084), .D(n6802), .Q(n7557) );
  OAI222 U1113 ( .A(n5060), .B(n10911), .C(n5036), .D(n6804), .Q(n7556) );
  OAI222 U1114 ( .A(n5012), .B(n10909), .C(n4988), .D(n6806), .Q(n7555) );
  OAI222 U1116 ( .A(n5348), .B(n10907), .C(n5324), .D(n6812), .Q(n7562) );
  OAI222 U1117 ( .A(n5300), .B(n10905), .C(n5276), .D(n6814), .Q(n7561) );
  OAI222 U1118 ( .A(n5252), .B(n10903), .C(n5228), .D(n6816), .Q(n7560) );
  OAI222 U1119 ( .A(n5204), .B(n10901), .C(n5180), .D(n6818), .Q(n7559) );
  OAI222 U1122 ( .A(n4004), .B(n10899), .C(n3980), .D(n6828), .Q(n7570) );
  OAI222 U1123 ( .A(n3956), .B(n10897), .C(n3932), .D(n6830), .Q(n7569) );
  OAI222 U1124 ( .A(n3908), .B(n10895), .C(n3884), .D(n6832), .Q(n7568) );
  OAI222 U1125 ( .A(n3860), .B(n10893), .C(n3836), .D(n6834), .Q(n7567) );
  OAI222 U1127 ( .A(n4196), .B(n10891), .C(n4172), .D(n6840), .Q(n7574) );
  OAI222 U1128 ( .A(n4148), .B(n10889), .C(n4124), .D(n6842), .Q(n7573) );
  OAI222 U1129 ( .A(n4100), .B(n10887), .C(n4076), .D(n6844), .Q(n7572) );
  OAI222 U1130 ( .A(n4052), .B(n10885), .C(n4028), .D(n6846), .Q(n7571) );
  OAI222 U1132 ( .A(n4388), .B(n10883), .C(n4364), .D(n6852), .Q(n7578) );
  OAI222 U1133 ( .A(n4340), .B(n10881), .C(n4316), .D(n6854), .Q(n7577) );
  OAI222 U1134 ( .A(n4292), .B(n6191), .C(n4268), .D(n6856), .Q(n7576) );
  OAI222 U1135 ( .A(n4244), .B(n6189), .C(n4220), .D(n6858), .Q(n7575) );
  OAI222 U1137 ( .A(n4580), .B(n6187), .C(n4556), .D(n6864), .Q(n7582) );
  OAI222 U1138 ( .A(n4532), .B(n6185), .C(n4508), .D(n6866), .Q(n7581) );
  OAI222 U1139 ( .A(n4484), .B(n6183), .C(n4460), .D(n6868), .Q(n7580) );
  OAI222 U1140 ( .A(n4436), .B(n6181), .C(n4412), .D(n6870), .Q(n7579) );
  OAI222 U1143 ( .A(n3236), .B(n6179), .C(n3212), .D(n6880), .Q(n7590) );
  OAI222 U1144 ( .A(n3188), .B(n6177), .C(n3164), .D(n6882), .Q(n7589) );
  OAI222 U1145 ( .A(n3140), .B(n6175), .C(n3116), .D(n6884), .Q(n7588) );
  OAI222 U1146 ( .A(n3092), .B(n6173), .C(n3068), .D(n6886), .Q(n7587) );
  OAI222 U1148 ( .A(n3428), .B(n6171), .C(n3404), .D(n6892), .Q(n7594) );
  OAI222 U1149 ( .A(n3380), .B(n6169), .C(n3356), .D(n6894), .Q(n7593) );
  OAI222 U1150 ( .A(n3332), .B(n6167), .C(n3308), .D(n6896), .Q(n7592) );
  OAI222 U1151 ( .A(n3284), .B(n6165), .C(n3260), .D(n6898), .Q(n7591) );
  OAI222 U1153 ( .A(n3620), .B(n6163), .C(n3596), .D(n6904), .Q(n7598) );
  OAI222 U1154 ( .A(n3572), .B(n6161), .C(n3548), .D(n6906), .Q(n7597) );
  OAI222 U1155 ( .A(n3524), .B(n6159), .C(n3500), .D(n6908), .Q(n7596) );
  OAI222 U1156 ( .A(n3476), .B(n6157), .C(n3452), .D(n6910), .Q(n7595) );
  OAI222 U1158 ( .A(n3812), .B(n6155), .C(n3788), .D(n6916), .Q(n7602) );
  OAI222 U1159 ( .A(n3764), .B(n6153), .C(n3740), .D(n6918), .Q(n7601) );
  OAI222 U1160 ( .A(n3716), .B(n6151), .C(n3692), .D(n6920), .Q(n7600) );
  OAI222 U1161 ( .A(n3668), .B(n6149), .C(n3644), .D(n6922), .Q(n7599) );
  OAI222 U1166 ( .A(n2467), .B(n11091), .C(n2443), .D(n6512), .Q(n7616) );
  OAI222 U1167 ( .A(n2419), .B(n11089), .C(n2395), .D(n6514), .Q(n7615) );
  OAI222 U1168 ( .A(n2371), .B(n11087), .C(n2347), .D(n6516), .Q(n7614) );
  OAI222 U1169 ( .A(n2323), .B(n11085), .C(n2299), .D(n6518), .Q(n7613) );
  OAI222 U1171 ( .A(n2659), .B(n11083), .C(n2635), .D(n6524), .Q(n7620) );
  OAI222 U1172 ( .A(n2611), .B(n11081), .C(n2587), .D(n6526), .Q(n7619) );
  OAI222 U1173 ( .A(n2563), .B(n11079), .C(n2539), .D(n6528), .Q(n7618) );
  OAI222 U1174 ( .A(n2515), .B(n11077), .C(n2491), .D(n6530), .Q(n7617) );
  OAI222 U1176 ( .A(n2851), .B(n11075), .C(n2827), .D(n6536), .Q(n7624) );
  OAI222 U1177 ( .A(n2803), .B(n11073), .C(n2779), .D(n6538), .Q(n7623) );
  OAI222 U1178 ( .A(n2755), .B(n11071), .C(n2731), .D(n6540), .Q(n7622) );
  OAI222 U1179 ( .A(n2707), .B(n11069), .C(n2683), .D(n6542), .Q(n7621) );
  OAI222 U1181 ( .A(n3043), .B(n11067), .C(n3019), .D(n6548), .Q(n7628) );
  OAI222 U1182 ( .A(n2995), .B(n11065), .C(n2971), .D(n6550), .Q(n7627) );
  OAI222 U1183 ( .A(n2947), .B(n11063), .C(n2923), .D(n6552), .Q(n7626) );
  OAI222 U1184 ( .A(n2899), .B(n11061), .C(n2875), .D(n6554), .Q(n7625) );
  OAI222 U1187 ( .A(n1699), .B(n11059), .C(n1675), .D(n6564), .Q(n7636) );
  OAI222 U1188 ( .A(n1651), .B(n11057), .C(n1627), .D(n6566), .Q(n7635) );
  OAI222 U1189 ( .A(n1603), .B(n11055), .C(n1579), .D(n6568), .Q(n7634) );
  OAI222 U1190 ( .A(n1555), .B(n11053), .C(n1531), .D(n6570), .Q(n7633) );
  OAI222 U1192 ( .A(n1891), .B(n11051), .C(n1867), .D(n6576), .Q(n7640) );
  OAI222 U1193 ( .A(n1843), .B(n11049), .C(n1819), .D(n6578), .Q(n7639) );
  OAI222 U1194 ( .A(n1795), .B(n11047), .C(n1771), .D(n6580), .Q(n7638) );
  OAI222 U1195 ( .A(n1747), .B(n11045), .C(n1723), .D(n6582), .Q(n7637) );
  OAI222 U1197 ( .A(n2083), .B(n11043), .C(n2059), .D(n6588), .Q(n7644) );
  OAI222 U1198 ( .A(n2035), .B(n11041), .C(n2011), .D(n6590), .Q(n7643) );
  OAI222 U1199 ( .A(n1987), .B(n11039), .C(n1963), .D(n6592), .Q(n7642) );
  OAI222 U1200 ( .A(n1939), .B(n11037), .C(n1915), .D(n6594), .Q(n7641) );
  OAI222 U1202 ( .A(n2275), .B(n11035), .C(n2251), .D(n6600), .Q(n7648) );
  OAI222 U1203 ( .A(n2227), .B(n11033), .C(n2203), .D(n6602), .Q(n7647) );
  OAI222 U1204 ( .A(n2179), .B(n11031), .C(n2155), .D(n6604), .Q(n7646) );
  OAI222 U1205 ( .A(n2131), .B(n11029), .C(n2107), .D(n6606), .Q(n7645) );
  OAI222 U1208 ( .A(n931), .B(n11027), .C(n907), .D(n6616), .Q(n7656) );
  OAI222 U1209 ( .A(n883), .B(n11025), .C(n859), .D(n6618), .Q(n7655) );
  OAI222 U1210 ( .A(n835), .B(n11023), .C(n811), .D(n6620), .Q(n7654) );
  OAI222 U1211 ( .A(n787), .B(n11021), .C(n763), .D(n6622), .Q(n7653) );
  OAI222 U1213 ( .A(n1123), .B(n11019), .C(n1099), .D(n6628), .Q(n7660) );
  OAI222 U1214 ( .A(n1075), .B(n11017), .C(n1051), .D(n6630), .Q(n7659) );
  OAI222 U1215 ( .A(n1027), .B(n11015), .C(n1003), .D(n6632), .Q(n7658) );
  OAI222 U1216 ( .A(n979), .B(n11013), .C(n955), .D(n6634), .Q(n7657) );
  OAI222 U1218 ( .A(n1315), .B(n11011), .C(n1291), .D(n6640), .Q(n7664) );
  OAI222 U1219 ( .A(n1267), .B(n11009), .C(n1243), .D(n6642), .Q(n7663) );
  OAI222 U1220 ( .A(n1219), .B(n11007), .C(n1195), .D(n6644), .Q(n7662) );
  OAI222 U1221 ( .A(n1171), .B(n11005), .C(n1147), .D(n6646), .Q(n7661) );
  OAI222 U1223 ( .A(n1507), .B(n11003), .C(n1483), .D(n6652), .Q(n7668) );
  OAI222 U1224 ( .A(n1459), .B(n11001), .C(n1435), .D(n6654), .Q(n7667) );
  OAI222 U1225 ( .A(n1411), .B(n10999), .C(n1387), .D(n6656), .Q(n7666) );
  OAI222 U1226 ( .A(n1363), .B(n10997), .C(n1339), .D(n6658), .Q(n7665) );
  OAI222 U1229 ( .A(n163), .B(n10995), .C(n139), .D(n6668), .Q(n7676) );
  OAI222 U1230 ( .A(n115), .B(n10993), .C(n91), .D(n6670), .Q(n7675) );
  OAI222 U1231 ( .A(n67), .B(n10991), .C(n43), .D(n6672), .Q(n7674) );
  OAI222 U1232 ( .A(n19), .B(n10989), .C(n6139), .D(n6674), .Q(n7673) );
  OAI222 U1234 ( .A(n355), .B(n10987), .C(n331), .D(n6680), .Q(n7680) );
  OAI222 U1235 ( .A(n307), .B(n10985), .C(n283), .D(n6682), .Q(n7679) );
  OAI222 U1236 ( .A(n259), .B(n10983), .C(n235), .D(n6684), .Q(n7678) );
  OAI222 U1237 ( .A(n211), .B(n10981), .C(n187), .D(n6686), .Q(n7677) );
  OAI222 U1239 ( .A(n547), .B(n10979), .C(n523), .D(n6692), .Q(n7684) );
  OAI222 U1240 ( .A(n499), .B(n10977), .C(n475), .D(n6694), .Q(n7683) );
  OAI222 U1241 ( .A(n451), .B(n10975), .C(n427), .D(n6696), .Q(n7682) );
  OAI222 U1242 ( .A(n403), .B(n10973), .C(n379), .D(n6698), .Q(n7681) );
  OAI222 U1244 ( .A(n739), .B(n10971), .C(n715), .D(n6704), .Q(n7688) );
  OAI222 U1245 ( .A(n691), .B(n10969), .C(n667), .D(n6706), .Q(n7687) );
  OAI222 U1246 ( .A(n643), .B(n10967), .C(n619), .D(n6708), .Q(n7686) );
  OAI222 U1247 ( .A(n595), .B(n10965), .C(n571), .D(n6710), .Q(n7685) );
  OAI222 U1251 ( .A(n5539), .B(n10963), .C(n5515), .D(n6724), .Q(n7700) );
  OAI222 U1252 ( .A(n5491), .B(n10961), .C(n5467), .D(n6726), .Q(n7699) );
  OAI222 U1253 ( .A(n5443), .B(n10959), .C(n5419), .D(n6728), .Q(n7698) );
  OAI222 U1254 ( .A(n5395), .B(n10957), .C(n5371), .D(n6730), .Q(n7697) );
  OAI222 U1256 ( .A(n5731), .B(n10955), .C(n5707), .D(n6736), .Q(n7704) );
  OAI222 U1257 ( .A(n5683), .B(n10953), .C(n5659), .D(n6738), .Q(n7703) );
  OAI222 U1258 ( .A(n5635), .B(n10951), .C(n5611), .D(n6740), .Q(n7702) );
  OAI222 U1259 ( .A(n5587), .B(n10949), .C(n5563), .D(n6742), .Q(n7701) );
  OAI222 U1261 ( .A(n5923), .B(n10947), .C(n5899), .D(n6748), .Q(n7708) );
  OAI222 U1262 ( .A(n5875), .B(n10945), .C(n5851), .D(n6750), .Q(n7707) );
  OAI222 U1263 ( .A(n5827), .B(n10943), .C(n5803), .D(n6752), .Q(n7706) );
  OAI222 U1264 ( .A(n5779), .B(n10941), .C(n5755), .D(n6754), .Q(n7705) );
  OAI222 U1266 ( .A(n6115), .B(n10939), .C(n6091), .D(n6760), .Q(n7712) );
  OAI222 U1267 ( .A(n6067), .B(n10937), .C(n6043), .D(n6762), .Q(n7711) );
  OAI222 U1268 ( .A(n6019), .B(n10935), .C(n5995), .D(n6764), .Q(n7710) );
  OAI222 U1269 ( .A(n5971), .B(n10933), .C(n5947), .D(n6766), .Q(n7709) );
  OAI222 U1272 ( .A(n4771), .B(n10931), .C(n4747), .D(n6776), .Q(n7720) );
  OAI222 U1273 ( .A(n4723), .B(n10929), .C(n4699), .D(n6778), .Q(n7719) );
  OAI222 U1274 ( .A(n4675), .B(n10927), .C(n4651), .D(n6780), .Q(n7718) );
  OAI222 U1275 ( .A(n4627), .B(n10925), .C(n4603), .D(n6782), .Q(n7717) );
  OAI222 U1277 ( .A(n4963), .B(n10923), .C(n4939), .D(n6788), .Q(n7724) );
  OAI222 U1278 ( .A(n4915), .B(n10921), .C(n4891), .D(n6790), .Q(n7723) );
  OAI222 U1279 ( .A(n4867), .B(n10919), .C(n4843), .D(n6792), .Q(n7722) );
  OAI222 U1280 ( .A(n4819), .B(n10917), .C(n4795), .D(n6794), .Q(n7721) );
  OAI222 U1282 ( .A(n5155), .B(n10915), .C(n5131), .D(n6800), .Q(n7728) );
  OAI222 U1283 ( .A(n5107), .B(n10913), .C(n5083), .D(n6802), .Q(n7727) );
  OAI222 U1284 ( .A(n5059), .B(n10911), .C(n5035), .D(n6804), .Q(n7726) );
  OAI222 U1285 ( .A(n5011), .B(n10909), .C(n4987), .D(n6806), .Q(n7725) );
  OAI222 U1287 ( .A(n5347), .B(n10907), .C(n5323), .D(n6812), .Q(n7732) );
  OAI222 U1288 ( .A(n5299), .B(n10905), .C(n5275), .D(n6814), .Q(n7731) );
  OAI222 U1289 ( .A(n5251), .B(n10903), .C(n5227), .D(n6816), .Q(n7730) );
  OAI222 U1290 ( .A(n5203), .B(n10901), .C(n5179), .D(n6818), .Q(n7729) );
  OAI222 U1293 ( .A(n4003), .B(n10899), .C(n3979), .D(n6828), .Q(n7740) );
  OAI222 U1294 ( .A(n3955), .B(n10897), .C(n3931), .D(n6830), .Q(n7739) );
  OAI222 U1295 ( .A(n3907), .B(n10895), .C(n3883), .D(n6832), .Q(n7738) );
  OAI222 U1296 ( .A(n3859), .B(n10893), .C(n3835), .D(n6834), .Q(n7737) );
  OAI222 U1298 ( .A(n4195), .B(n10891), .C(n4171), .D(n6840), .Q(n7744) );
  OAI222 U1299 ( .A(n4147), .B(n10889), .C(n4123), .D(n6842), .Q(n7743) );
  OAI222 U1300 ( .A(n4099), .B(n10887), .C(n4075), .D(n6844), .Q(n7742) );
  OAI222 U1301 ( .A(n4051), .B(n10885), .C(n4027), .D(n6846), .Q(n7741) );
  OAI222 U1303 ( .A(n4387), .B(n10883), .C(n4363), .D(n6852), .Q(n7748) );
  OAI222 U1304 ( .A(n4339), .B(n10881), .C(n4315), .D(n6854), .Q(n7747) );
  OAI222 U1305 ( .A(n4291), .B(n6191), .C(n4267), .D(n6856), .Q(n7746) );
  OAI222 U1306 ( .A(n4243), .B(n6189), .C(n4219), .D(n6858), .Q(n7745) );
  OAI222 U1308 ( .A(n4579), .B(n6187), .C(n4555), .D(n6864), .Q(n7752) );
  OAI222 U1309 ( .A(n4531), .B(n6185), .C(n4507), .D(n6866), .Q(n7751) );
  OAI222 U1310 ( .A(n4483), .B(n6183), .C(n4459), .D(n6868), .Q(n7750) );
  OAI222 U1311 ( .A(n4435), .B(n6181), .C(n4411), .D(n6870), .Q(n7749) );
  OAI222 U1314 ( .A(n3235), .B(n6179), .C(n3211), .D(n6880), .Q(n7760) );
  OAI222 U1315 ( .A(n3187), .B(n6177), .C(n3163), .D(n6882), .Q(n7759) );
  OAI222 U1316 ( .A(n3139), .B(n6175), .C(n3115), .D(n6884), .Q(n7758) );
  OAI222 U1317 ( .A(n3091), .B(n6173), .C(n3067), .D(n6886), .Q(n7757) );
  OAI222 U1319 ( .A(n3427), .B(n6171), .C(n3403), .D(n6892), .Q(n7764) );
  OAI222 U1320 ( .A(n3379), .B(n6169), .C(n3355), .D(n6894), .Q(n7763) );
  OAI222 U1321 ( .A(n3331), .B(n6167), .C(n3307), .D(n6896), .Q(n7762) );
  OAI222 U1322 ( .A(n3283), .B(n6165), .C(n3259), .D(n6898), .Q(n7761) );
  OAI222 U1324 ( .A(n3619), .B(n6163), .C(n3595), .D(n6904), .Q(n7768) );
  OAI222 U1325 ( .A(n3571), .B(n6161), .C(n3547), .D(n6906), .Q(n7767) );
  OAI222 U1326 ( .A(n3523), .B(n6159), .C(n3499), .D(n6908), .Q(n7766) );
  OAI222 U1327 ( .A(n3475), .B(n6157), .C(n3451), .D(n6910), .Q(n7765) );
  OAI222 U1329 ( .A(n3811), .B(n6155), .C(n3787), .D(n6916), .Q(n7772) );
  OAI222 U1330 ( .A(n3763), .B(n6153), .C(n3739), .D(n6918), .Q(n7771) );
  OAI222 U1331 ( .A(n3715), .B(n6151), .C(n3691), .D(n6920), .Q(n7770) );
  OAI222 U1332 ( .A(n3667), .B(n6149), .C(n3643), .D(n6922), .Q(n7769) );
  OAI222 U1337 ( .A(n2466), .B(n11091), .C(n2442), .D(n6512), .Q(n7786) );
  OAI222 U1338 ( .A(n2418), .B(n11089), .C(n2394), .D(n6514), .Q(n7785) );
  OAI222 U1339 ( .A(n2370), .B(n11087), .C(n2346), .D(n6516), .Q(n7784) );
  OAI222 U1340 ( .A(n2322), .B(n11085), .C(n2298), .D(n6518), .Q(n7783) );
  OAI222 U1342 ( .A(n2658), .B(n11083), .C(n2634), .D(n6524), .Q(n7790) );
  OAI222 U1343 ( .A(n2610), .B(n11081), .C(n2586), .D(n6526), .Q(n7789) );
  OAI222 U1344 ( .A(n2562), .B(n11079), .C(n2538), .D(n6528), .Q(n7788) );
  OAI222 U1345 ( .A(n2514), .B(n11077), .C(n2490), .D(n6530), .Q(n7787) );
  OAI222 U1347 ( .A(n2850), .B(n11075), .C(n2826), .D(n6536), .Q(n7794) );
  OAI222 U1348 ( .A(n2802), .B(n11073), .C(n2778), .D(n6538), .Q(n7793) );
  OAI222 U1349 ( .A(n2754), .B(n11071), .C(n2730), .D(n6540), .Q(n7792) );
  OAI222 U1350 ( .A(n2706), .B(n11069), .C(n2682), .D(n6542), .Q(n7791) );
  OAI222 U1352 ( .A(n3042), .B(n11067), .C(n3018), .D(n6548), .Q(n7798) );
  OAI222 U1353 ( .A(n2994), .B(n11065), .C(n2970), .D(n6550), .Q(n7797) );
  OAI222 U1354 ( .A(n2946), .B(n11063), .C(n2922), .D(n6552), .Q(n7796) );
  OAI222 U1355 ( .A(n2898), .B(n11061), .C(n2874), .D(n6554), .Q(n7795) );
  OAI222 U1358 ( .A(n1698), .B(n11059), .C(n1674), .D(n6564), .Q(n7806) );
  OAI222 U1359 ( .A(n1650), .B(n11057), .C(n1626), .D(n6566), .Q(n7805) );
  OAI222 U1360 ( .A(n1602), .B(n11055), .C(n1578), .D(n6568), .Q(n7804) );
  OAI222 U1361 ( .A(n1554), .B(n11053), .C(n1530), .D(n6570), .Q(n7803) );
  OAI222 U1363 ( .A(n1890), .B(n11051), .C(n1866), .D(n6576), .Q(n7810) );
  OAI222 U1364 ( .A(n1842), .B(n11049), .C(n1818), .D(n6578), .Q(n7809) );
  OAI222 U1365 ( .A(n1794), .B(n11047), .C(n1770), .D(n6580), .Q(n7808) );
  OAI222 U1366 ( .A(n1746), .B(n11045), .C(n1722), .D(n6582), .Q(n7807) );
  OAI222 U1368 ( .A(n2082), .B(n11043), .C(n2058), .D(n6588), .Q(n7814) );
  OAI222 U1369 ( .A(n2034), .B(n11041), .C(n2010), .D(n6590), .Q(n7813) );
  OAI222 U1370 ( .A(n1986), .B(n11039), .C(n1962), .D(n6592), .Q(n7812) );
  OAI222 U1371 ( .A(n1938), .B(n11037), .C(n1914), .D(n6594), .Q(n7811) );
  OAI222 U1373 ( .A(n2274), .B(n11035), .C(n2250), .D(n6600), .Q(n7818) );
  OAI222 U1374 ( .A(n2226), .B(n11033), .C(n2202), .D(n6602), .Q(n7817) );
  OAI222 U1375 ( .A(n2178), .B(n11031), .C(n2154), .D(n6604), .Q(n7816) );
  OAI222 U1376 ( .A(n2130), .B(n11029), .C(n2106), .D(n6606), .Q(n7815) );
  OAI222 U1379 ( .A(n930), .B(n11027), .C(n906), .D(n6616), .Q(n7826) );
  OAI222 U1380 ( .A(n882), .B(n11025), .C(n858), .D(n6618), .Q(n7825) );
  OAI222 U1381 ( .A(n834), .B(n11023), .C(n810), .D(n6620), .Q(n7824) );
  OAI222 U1382 ( .A(n786), .B(n11021), .C(n762), .D(n6622), .Q(n7823) );
  OAI222 U1384 ( .A(n1122), .B(n11019), .C(n1098), .D(n6628), .Q(n7830) );
  OAI222 U1385 ( .A(n1074), .B(n11017), .C(n1050), .D(n6630), .Q(n7829) );
  OAI222 U1386 ( .A(n1026), .B(n11015), .C(n1002), .D(n6632), .Q(n7828) );
  OAI222 U1387 ( .A(n978), .B(n11013), .C(n954), .D(n6634), .Q(n7827) );
  OAI222 U1389 ( .A(n1314), .B(n11011), .C(n1290), .D(n6640), .Q(n7834) );
  OAI222 U1390 ( .A(n1266), .B(n11009), .C(n1242), .D(n6642), .Q(n7833) );
  OAI222 U1391 ( .A(n1218), .B(n11007), .C(n1194), .D(n6644), .Q(n7832) );
  OAI222 U1392 ( .A(n1170), .B(n11005), .C(n1146), .D(n6646), .Q(n7831) );
  OAI222 U1394 ( .A(n1506), .B(n11003), .C(n1482), .D(n6652), .Q(n7838) );
  OAI222 U1395 ( .A(n1458), .B(n11001), .C(n1434), .D(n6654), .Q(n7837) );
  OAI222 U1396 ( .A(n1410), .B(n10999), .C(n1386), .D(n6656), .Q(n7836) );
  OAI222 U1397 ( .A(n1362), .B(n10997), .C(n1338), .D(n6658), .Q(n7835) );
  OAI222 U1400 ( .A(n162), .B(n10995), .C(n138), .D(n6668), .Q(n7846) );
  OAI222 U1401 ( .A(n114), .B(n10993), .C(n90), .D(n6670), .Q(n7845) );
  OAI222 U1402 ( .A(n66), .B(n10991), .C(n42), .D(n6672), .Q(n7844) );
  OAI222 U1403 ( .A(n18), .B(n10989), .C(n6138), .D(n6674), .Q(n7843) );
  OAI222 U1405 ( .A(n354), .B(n10987), .C(n330), .D(n6680), .Q(n7850) );
  OAI222 U1406 ( .A(n306), .B(n10985), .C(n282), .D(n6682), .Q(n7849) );
  OAI222 U1407 ( .A(n258), .B(n10983), .C(n234), .D(n6684), .Q(n7848) );
  OAI222 U1408 ( .A(n210), .B(n10981), .C(n186), .D(n6686), .Q(n7847) );
  OAI222 U1410 ( .A(n546), .B(n10979), .C(n522), .D(n6692), .Q(n7854) );
  OAI222 U1411 ( .A(n498), .B(n10977), .C(n474), .D(n6694), .Q(n7853) );
  OAI222 U1412 ( .A(n450), .B(n10975), .C(n426), .D(n6696), .Q(n7852) );
  OAI222 U1413 ( .A(n402), .B(n10973), .C(n378), .D(n6698), .Q(n7851) );
  OAI222 U1415 ( .A(n738), .B(n10971), .C(n714), .D(n6704), .Q(n7858) );
  OAI222 U1416 ( .A(n690), .B(n10969), .C(n666), .D(n6706), .Q(n7857) );
  OAI222 U1417 ( .A(n642), .B(n10967), .C(n618), .D(n6708), .Q(n7856) );
  OAI222 U1418 ( .A(n594), .B(n10965), .C(n570), .D(n6710), .Q(n7855) );
  OAI222 U1422 ( .A(n5538), .B(n10963), .C(n5514), .D(n6724), .Q(n7870) );
  OAI222 U1423 ( .A(n5490), .B(n10961), .C(n5466), .D(n6726), .Q(n7869) );
  OAI222 U1424 ( .A(n5442), .B(n10959), .C(n5418), .D(n6728), .Q(n7868) );
  OAI222 U1425 ( .A(n5394), .B(n10957), .C(n5370), .D(n6730), .Q(n7867) );
  OAI222 U1427 ( .A(n5730), .B(n10955), .C(n5706), .D(n6736), .Q(n7874) );
  OAI222 U1428 ( .A(n5682), .B(n10953), .C(n5658), .D(n6738), .Q(n7873) );
  OAI222 U1429 ( .A(n5634), .B(n10951), .C(n5610), .D(n6740), .Q(n7872) );
  OAI222 U1430 ( .A(n5586), .B(n10949), .C(n5562), .D(n6742), .Q(n7871) );
  OAI222 U1432 ( .A(n5922), .B(n10947), .C(n5898), .D(n6748), .Q(n7878) );
  OAI222 U1433 ( .A(n5874), .B(n10945), .C(n5850), .D(n6750), .Q(n7877) );
  OAI222 U1434 ( .A(n5826), .B(n10943), .C(n5802), .D(n6752), .Q(n7876) );
  OAI222 U1435 ( .A(n5778), .B(n10941), .C(n5754), .D(n6754), .Q(n7875) );
  OAI222 U1437 ( .A(n6114), .B(n10939), .C(n6090), .D(n6760), .Q(n7882) );
  OAI222 U1438 ( .A(n6066), .B(n10937), .C(n6042), .D(n6762), .Q(n7881) );
  OAI222 U1439 ( .A(n6018), .B(n10935), .C(n5994), .D(n6764), .Q(n7880) );
  OAI222 U1440 ( .A(n5970), .B(n10933), .C(n5946), .D(n6766), .Q(n7879) );
  OAI222 U1443 ( .A(n4770), .B(n10931), .C(n4746), .D(n6776), .Q(n7890) );
  OAI222 U1444 ( .A(n4722), .B(n10929), .C(n4698), .D(n6778), .Q(n7889) );
  OAI222 U1445 ( .A(n4674), .B(n10927), .C(n4650), .D(n6780), .Q(n7888) );
  OAI222 U1446 ( .A(n4626), .B(n10925), .C(n4602), .D(n6782), .Q(n7887) );
  OAI222 U1448 ( .A(n4962), .B(n10923), .C(n4938), .D(n6788), .Q(n7894) );
  OAI222 U1449 ( .A(n4914), .B(n10921), .C(n4890), .D(n6790), .Q(n7893) );
  OAI222 U1450 ( .A(n4866), .B(n10919), .C(n4842), .D(n6792), .Q(n7892) );
  OAI222 U1451 ( .A(n4818), .B(n10917), .C(n4794), .D(n6794), .Q(n7891) );
  OAI222 U1453 ( .A(n5154), .B(n10915), .C(n5130), .D(n6800), .Q(n7898) );
  OAI222 U1454 ( .A(n5106), .B(n10913), .C(n5082), .D(n6802), .Q(n7897) );
  OAI222 U1455 ( .A(n5058), .B(n10911), .C(n5034), .D(n6804), .Q(n7896) );
  OAI222 U1456 ( .A(n5010), .B(n10909), .C(n4986), .D(n6806), .Q(n7895) );
  OAI222 U1458 ( .A(n5346), .B(n10907), .C(n5322), .D(n6812), .Q(n7902) );
  OAI222 U1459 ( .A(n5298), .B(n10905), .C(n5274), .D(n6814), .Q(n7901) );
  OAI222 U1460 ( .A(n5250), .B(n10903), .C(n5226), .D(n6816), .Q(n7900) );
  OAI222 U1461 ( .A(n5202), .B(n10901), .C(n5178), .D(n6818), .Q(n7899) );
  OAI222 U1464 ( .A(n4002), .B(n10899), .C(n3978), .D(n6828), .Q(n7910) );
  OAI222 U1465 ( .A(n3954), .B(n10897), .C(n3930), .D(n6830), .Q(n7909) );
  OAI222 U1466 ( .A(n3906), .B(n10895), .C(n3882), .D(n6832), .Q(n7908) );
  OAI222 U1467 ( .A(n3858), .B(n10893), .C(n3834), .D(n6834), .Q(n7907) );
  OAI222 U1469 ( .A(n4194), .B(n10891), .C(n4170), .D(n6840), .Q(n7914) );
  OAI222 U1470 ( .A(n4146), .B(n10889), .C(n4122), .D(n6842), .Q(n7913) );
  OAI222 U1471 ( .A(n4098), .B(n10887), .C(n4074), .D(n6844), .Q(n7912) );
  OAI222 U1472 ( .A(n4050), .B(n10885), .C(n4026), .D(n6846), .Q(n7911) );
  OAI222 U1474 ( .A(n4386), .B(n10883), .C(n4362), .D(n6852), .Q(n7918) );
  OAI222 U1475 ( .A(n4338), .B(n10881), .C(n4314), .D(n6854), .Q(n7917) );
  OAI222 U1476 ( .A(n4290), .B(n6191), .C(n4266), .D(n6856), .Q(n7916) );
  OAI222 U1477 ( .A(n4242), .B(n6189), .C(n4218), .D(n6858), .Q(n7915) );
  OAI222 U1479 ( .A(n4578), .B(n6187), .C(n4554), .D(n6864), .Q(n7922) );
  OAI222 U1480 ( .A(n4530), .B(n6185), .C(n4506), .D(n6866), .Q(n7921) );
  OAI222 U1481 ( .A(n4482), .B(n6183), .C(n4458), .D(n6868), .Q(n7920) );
  OAI222 U1482 ( .A(n4434), .B(n6181), .C(n4410), .D(n6870), .Q(n7919) );
  OAI222 U1485 ( .A(n3234), .B(n6179), .C(n3210), .D(n6880), .Q(n7930) );
  OAI222 U1486 ( .A(n3186), .B(n6177), .C(n3162), .D(n6882), .Q(n7929) );
  OAI222 U1487 ( .A(n3138), .B(n6175), .C(n3114), .D(n6884), .Q(n7928) );
  OAI222 U1488 ( .A(n3090), .B(n6173), .C(n3066), .D(n6886), .Q(n7927) );
  OAI222 U1490 ( .A(n3426), .B(n6171), .C(n3402), .D(n6892), .Q(n7934) );
  OAI222 U1491 ( .A(n3378), .B(n6169), .C(n3354), .D(n6894), .Q(n7933) );
  OAI222 U1492 ( .A(n3330), .B(n6167), .C(n3306), .D(n6896), .Q(n7932) );
  OAI222 U1493 ( .A(n3282), .B(n6165), .C(n3258), .D(n6898), .Q(n7931) );
  OAI222 U1495 ( .A(n3618), .B(n6163), .C(n3594), .D(n6904), .Q(n7938) );
  OAI222 U1496 ( .A(n3570), .B(n6161), .C(n3546), .D(n6906), .Q(n7937) );
  OAI222 U1497 ( .A(n3522), .B(n6159), .C(n3498), .D(n6908), .Q(n7936) );
  OAI222 U1498 ( .A(n3474), .B(n6157), .C(n3450), .D(n6910), .Q(n7935) );
  OAI222 U1500 ( .A(n3810), .B(n6155), .C(n3786), .D(n6916), .Q(n7942) );
  OAI222 U1501 ( .A(n3762), .B(n6153), .C(n3738), .D(n6918), .Q(n7941) );
  OAI222 U1502 ( .A(n3714), .B(n6151), .C(n3690), .D(n6920), .Q(n7940) );
  OAI222 U1503 ( .A(n3666), .B(n6149), .C(n3642), .D(n6922), .Q(n7939) );
  OAI222 U1508 ( .A(n2465), .B(n11091), .C(n2441), .D(n6512), .Q(n7956) );
  OAI222 U1509 ( .A(n2417), .B(n11089), .C(n2393), .D(n6514), .Q(n7955) );
  OAI222 U1510 ( .A(n2369), .B(n11087), .C(n2345), .D(n6516), .Q(n7954) );
  OAI222 U1511 ( .A(n2321), .B(n11085), .C(n2297), .D(n6518), .Q(n7953) );
  OAI222 U1513 ( .A(n2657), .B(n11083), .C(n2633), .D(n6524), .Q(n7960) );
  OAI222 U1514 ( .A(n2609), .B(n11081), .C(n2585), .D(n6526), .Q(n7959) );
  OAI222 U1515 ( .A(n2561), .B(n11079), .C(n2537), .D(n6528), .Q(n7958) );
  OAI222 U1516 ( .A(n2513), .B(n11077), .C(n2489), .D(n6530), .Q(n7957) );
  OAI222 U1518 ( .A(n2849), .B(n11075), .C(n2825), .D(n6536), .Q(n7964) );
  OAI222 U1519 ( .A(n2801), .B(n11073), .C(n2777), .D(n6538), .Q(n7963) );
  OAI222 U1520 ( .A(n2753), .B(n11071), .C(n2729), .D(n6540), .Q(n7962) );
  OAI222 U1521 ( .A(n2705), .B(n11069), .C(n2681), .D(n6542), .Q(n7961) );
  OAI222 U1523 ( .A(n3041), .B(n11067), .C(n3017), .D(n6548), .Q(n7968) );
  OAI222 U1524 ( .A(n2993), .B(n11065), .C(n2969), .D(n6550), .Q(n7967) );
  OAI222 U1525 ( .A(n2945), .B(n11063), .C(n2921), .D(n6552), .Q(n7966) );
  OAI222 U1526 ( .A(n2897), .B(n11061), .C(n2873), .D(n6554), .Q(n7965) );
  OAI222 U1529 ( .A(n1697), .B(n11059), .C(n1673), .D(n6564), .Q(n7976) );
  OAI222 U1530 ( .A(n1649), .B(n11057), .C(n1625), .D(n6566), .Q(n7975) );
  OAI222 U1531 ( .A(n1601), .B(n11055), .C(n1577), .D(n6568), .Q(n7974) );
  OAI222 U1532 ( .A(n1553), .B(n11053), .C(n1529), .D(n6570), .Q(n7973) );
  OAI222 U1534 ( .A(n1889), .B(n11051), .C(n1865), .D(n6576), .Q(n7980) );
  OAI222 U1535 ( .A(n1841), .B(n11049), .C(n1817), .D(n6578), .Q(n7979) );
  OAI222 U1536 ( .A(n1793), .B(n11047), .C(n1769), .D(n6580), .Q(n7978) );
  OAI222 U1537 ( .A(n1745), .B(n11045), .C(n1721), .D(n6582), .Q(n7977) );
  OAI222 U1539 ( .A(n2081), .B(n11043), .C(n2057), .D(n6588), .Q(n7984) );
  OAI222 U1540 ( .A(n2033), .B(n11041), .C(n2009), .D(n6590), .Q(n7983) );
  OAI222 U1541 ( .A(n1985), .B(n11039), .C(n1961), .D(n6592), .Q(n7982) );
  OAI222 U1542 ( .A(n1937), .B(n11037), .C(n1913), .D(n6594), .Q(n7981) );
  OAI222 U1544 ( .A(n2273), .B(n11035), .C(n2249), .D(n6600), .Q(n7988) );
  OAI222 U1545 ( .A(n2225), .B(n11033), .C(n2201), .D(n6602), .Q(n7987) );
  OAI222 U1546 ( .A(n2177), .B(n11031), .C(n2153), .D(n6604), .Q(n7986) );
  OAI222 U1547 ( .A(n2129), .B(n11029), .C(n2105), .D(n6606), .Q(n7985) );
  OAI222 U1550 ( .A(n929), .B(n11027), .C(n905), .D(n6616), .Q(n7996) );
  OAI222 U1551 ( .A(n881), .B(n11025), .C(n857), .D(n6618), .Q(n7995) );
  OAI222 U1552 ( .A(n833), .B(n11023), .C(n809), .D(n6620), .Q(n7994) );
  OAI222 U1553 ( .A(n785), .B(n11021), .C(n761), .D(n6622), .Q(n7993) );
  OAI222 U1555 ( .A(n1121), .B(n11019), .C(n1097), .D(n6628), .Q(n8000) );
  OAI222 U1556 ( .A(n1073), .B(n11017), .C(n1049), .D(n6630), .Q(n7999) );
  OAI222 U1557 ( .A(n1025), .B(n11015), .C(n1001), .D(n6632), .Q(n7998) );
  OAI222 U1558 ( .A(n977), .B(n11013), .C(n953), .D(n6634), .Q(n7997) );
  OAI222 U1560 ( .A(n1313), .B(n11011), .C(n1289), .D(n6640), .Q(n8004) );
  OAI222 U1561 ( .A(n1265), .B(n11009), .C(n1241), .D(n6642), .Q(n8003) );
  OAI222 U1562 ( .A(n1217), .B(n11007), .C(n1193), .D(n6644), .Q(n8002) );
  OAI222 U1563 ( .A(n1169), .B(n11005), .C(n1145), .D(n6646), .Q(n8001) );
  OAI222 U1565 ( .A(n1505), .B(n11003), .C(n1481), .D(n6652), .Q(n8008) );
  OAI222 U1566 ( .A(n1457), .B(n11001), .C(n1433), .D(n6654), .Q(n8007) );
  OAI222 U1567 ( .A(n1409), .B(n10999), .C(n1385), .D(n6656), .Q(n8006) );
  OAI222 U1568 ( .A(n1361), .B(n10997), .C(n1337), .D(n6658), .Q(n8005) );
  OAI222 U1571 ( .A(n161), .B(n10995), .C(n137), .D(n6668), .Q(n8016) );
  OAI222 U1572 ( .A(n113), .B(n10993), .C(n89), .D(n6670), .Q(n8015) );
  OAI222 U1573 ( .A(n65), .B(n10991), .C(n41), .D(n6672), .Q(n8014) );
  OAI222 U1574 ( .A(n17), .B(n10989), .C(n6137), .D(n6674), .Q(n8013) );
  OAI222 U1576 ( .A(n353), .B(n10987), .C(n329), .D(n6680), .Q(n8020) );
  OAI222 U1577 ( .A(n305), .B(n10985), .C(n281), .D(n6682), .Q(n8019) );
  OAI222 U1578 ( .A(n257), .B(n10983), .C(n233), .D(n6684), .Q(n8018) );
  OAI222 U1579 ( .A(n209), .B(n10981), .C(n185), .D(n6686), .Q(n8017) );
  OAI222 U1581 ( .A(n545), .B(n10979), .C(n521), .D(n6692), .Q(n8024) );
  OAI222 U1582 ( .A(n497), .B(n10977), .C(n473), .D(n6694), .Q(n8023) );
  OAI222 U1583 ( .A(n449), .B(n10975), .C(n425), .D(n6696), .Q(n8022) );
  OAI222 U1584 ( .A(n401), .B(n10973), .C(n377), .D(n6698), .Q(n8021) );
  OAI222 U1586 ( .A(n737), .B(n10971), .C(n713), .D(n6704), .Q(n8028) );
  OAI222 U1587 ( .A(n689), .B(n10969), .C(n665), .D(n6706), .Q(n8027) );
  OAI222 U1588 ( .A(n641), .B(n10967), .C(n617), .D(n6708), .Q(n8026) );
  OAI222 U1589 ( .A(n593), .B(n10965), .C(n569), .D(n6710), .Q(n8025) );
  OAI222 U1593 ( .A(n5537), .B(n10963), .C(n5513), .D(n6724), .Q(n8040) );
  OAI222 U1594 ( .A(n5489), .B(n10961), .C(n5465), .D(n6726), .Q(n8039) );
  OAI222 U1595 ( .A(n5441), .B(n10959), .C(n5417), .D(n6728), .Q(n8038) );
  OAI222 U1596 ( .A(n5393), .B(n10957), .C(n5369), .D(n6730), .Q(n8037) );
  OAI222 U1598 ( .A(n5729), .B(n10955), .C(n5705), .D(n6736), .Q(n8044) );
  OAI222 U1599 ( .A(n5681), .B(n10953), .C(n5657), .D(n6738), .Q(n8043) );
  OAI222 U1600 ( .A(n5633), .B(n10951), .C(n5609), .D(n6740), .Q(n8042) );
  OAI222 U1601 ( .A(n5585), .B(n10949), .C(n5561), .D(n6742), .Q(n8041) );
  OAI222 U1603 ( .A(n5921), .B(n10947), .C(n5897), .D(n6748), .Q(n8048) );
  OAI222 U1604 ( .A(n5873), .B(n10945), .C(n5849), .D(n6750), .Q(n8047) );
  OAI222 U1605 ( .A(n5825), .B(n10943), .C(n5801), .D(n6752), .Q(n8046) );
  OAI222 U1606 ( .A(n5777), .B(n10941), .C(n5753), .D(n6754), .Q(n8045) );
  OAI222 U1608 ( .A(n6113), .B(n10939), .C(n6089), .D(n6760), .Q(n8052) );
  OAI222 U1609 ( .A(n6065), .B(n10937), .C(n6041), .D(n6762), .Q(n8051) );
  OAI222 U1610 ( .A(n6017), .B(n10935), .C(n5993), .D(n6764), .Q(n8050) );
  OAI222 U1611 ( .A(n5969), .B(n10933), .C(n5945), .D(n6766), .Q(n8049) );
  OAI222 U1614 ( .A(n4769), .B(n10931), .C(n4745), .D(n6776), .Q(n8060) );
  OAI222 U1615 ( .A(n4721), .B(n10929), .C(n4697), .D(n6778), .Q(n8059) );
  OAI222 U1616 ( .A(n4673), .B(n10927), .C(n4649), .D(n6780), .Q(n8058) );
  OAI222 U1617 ( .A(n4625), .B(n10925), .C(n4601), .D(n6782), .Q(n8057) );
  OAI222 U1619 ( .A(n4961), .B(n10923), .C(n4937), .D(n6788), .Q(n8064) );
  OAI222 U1620 ( .A(n4913), .B(n10921), .C(n4889), .D(n6790), .Q(n8063) );
  OAI222 U1621 ( .A(n4865), .B(n10919), .C(n4841), .D(n6792), .Q(n8062) );
  OAI222 U1622 ( .A(n4817), .B(n10917), .C(n4793), .D(n6794), .Q(n8061) );
  OAI222 U1624 ( .A(n5153), .B(n10915), .C(n5129), .D(n6800), .Q(n8068) );
  OAI222 U1625 ( .A(n5105), .B(n10913), .C(n5081), .D(n6802), .Q(n8067) );
  OAI222 U1626 ( .A(n5057), .B(n10911), .C(n5033), .D(n6804), .Q(n8066) );
  OAI222 U1627 ( .A(n5009), .B(n10909), .C(n4985), .D(n6806), .Q(n8065) );
  OAI222 U1629 ( .A(n5345), .B(n10907), .C(n5321), .D(n6812), .Q(n8072) );
  OAI222 U1630 ( .A(n5297), .B(n10905), .C(n5273), .D(n6814), .Q(n8071) );
  OAI222 U1631 ( .A(n5249), .B(n10903), .C(n5225), .D(n6816), .Q(n8070) );
  OAI222 U1632 ( .A(n5201), .B(n10901), .C(n5177), .D(n6818), .Q(n8069) );
  OAI222 U1635 ( .A(n4001), .B(n10899), .C(n3977), .D(n6828), .Q(n8080) );
  OAI222 U1636 ( .A(n3953), .B(n10897), .C(n3929), .D(n6830), .Q(n8079) );
  OAI222 U1637 ( .A(n3905), .B(n10895), .C(n3881), .D(n6832), .Q(n8078) );
  OAI222 U1638 ( .A(n3857), .B(n10893), .C(n3833), .D(n6834), .Q(n8077) );
  OAI222 U1640 ( .A(n4193), .B(n10891), .C(n4169), .D(n6840), .Q(n8084) );
  OAI222 U1641 ( .A(n4145), .B(n10889), .C(n4121), .D(n6842), .Q(n8083) );
  OAI222 U1642 ( .A(n4097), .B(n10887), .C(n4073), .D(n6844), .Q(n8082) );
  OAI222 U1643 ( .A(n4049), .B(n10885), .C(n4025), .D(n6846), .Q(n8081) );
  OAI222 U1645 ( .A(n4385), .B(n10883), .C(n4361), .D(n6852), .Q(n8088) );
  OAI222 U1646 ( .A(n4337), .B(n10881), .C(n4313), .D(n6854), .Q(n8087) );
  OAI222 U1647 ( .A(n4289), .B(n6191), .C(n4265), .D(n6856), .Q(n8086) );
  OAI222 U1648 ( .A(n4241), .B(n6189), .C(n4217), .D(n6858), .Q(n8085) );
  OAI222 U1650 ( .A(n4577), .B(n6187), .C(n4553), .D(n6864), .Q(n8092) );
  OAI222 U1651 ( .A(n4529), .B(n6185), .C(n4505), .D(n6866), .Q(n8091) );
  OAI222 U1652 ( .A(n4481), .B(n6183), .C(n4457), .D(n6868), .Q(n8090) );
  OAI222 U1653 ( .A(n4433), .B(n6181), .C(n4409), .D(n6870), .Q(n8089) );
  OAI222 U1656 ( .A(n3233), .B(n6179), .C(n3209), .D(n6880), .Q(n8100) );
  OAI222 U1657 ( .A(n3185), .B(n6177), .C(n3161), .D(n6882), .Q(n8099) );
  OAI222 U1658 ( .A(n3137), .B(n6175), .C(n3113), .D(n6884), .Q(n8098) );
  OAI222 U1659 ( .A(n3089), .B(n6173), .C(n3065), .D(n6886), .Q(n8097) );
  OAI222 U1661 ( .A(n3425), .B(n6171), .C(n3401), .D(n6892), .Q(n8104) );
  OAI222 U1662 ( .A(n3377), .B(n6169), .C(n3353), .D(n6894), .Q(n8103) );
  OAI222 U1663 ( .A(n3329), .B(n6167), .C(n3305), .D(n6896), .Q(n8102) );
  OAI222 U1664 ( .A(n3281), .B(n6165), .C(n3257), .D(n6898), .Q(n8101) );
  OAI222 U1666 ( .A(n3617), .B(n6163), .C(n3593), .D(n6904), .Q(n8108) );
  OAI222 U1667 ( .A(n3569), .B(n6161), .C(n3545), .D(n6906), .Q(n8107) );
  OAI222 U1668 ( .A(n3521), .B(n6159), .C(n3497), .D(n6908), .Q(n8106) );
  OAI222 U1669 ( .A(n3473), .B(n6157), .C(n3449), .D(n6910), .Q(n8105) );
  OAI222 U1671 ( .A(n3809), .B(n6155), .C(n3785), .D(n6916), .Q(n8112) );
  OAI222 U1672 ( .A(n3761), .B(n6153), .C(n3737), .D(n6918), .Q(n8111) );
  OAI222 U1673 ( .A(n3713), .B(n6151), .C(n3689), .D(n6920), .Q(n8110) );
  OAI222 U1674 ( .A(n3665), .B(n6149), .C(n3641), .D(n6922), .Q(n8109) );
  OAI222 U1679 ( .A(n2464), .B(n11091), .C(n2440), .D(n6512), .Q(n8126) );
  OAI222 U1680 ( .A(n2416), .B(n11089), .C(n2392), .D(n6514), .Q(n8125) );
  OAI222 U1681 ( .A(n2368), .B(n11087), .C(n2344), .D(n6516), .Q(n8124) );
  OAI222 U1682 ( .A(n2320), .B(n11085), .C(n2296), .D(n6518), .Q(n8123) );
  OAI222 U1684 ( .A(n2656), .B(n11083), .C(n2632), .D(n6524), .Q(n8130) );
  OAI222 U1685 ( .A(n2608), .B(n11081), .C(n2584), .D(n6526), .Q(n8129) );
  OAI222 U1686 ( .A(n2560), .B(n11079), .C(n2536), .D(n6528), .Q(n8128) );
  OAI222 U1687 ( .A(n2512), .B(n11077), .C(n2488), .D(n6530), .Q(n8127) );
  OAI222 U1689 ( .A(n2848), .B(n11075), .C(n2824), .D(n6536), .Q(n8134) );
  OAI222 U1690 ( .A(n2800), .B(n11073), .C(n2776), .D(n6538), .Q(n8133) );
  OAI222 U1691 ( .A(n2752), .B(n11071), .C(n2728), .D(n6540), .Q(n8132) );
  OAI222 U1692 ( .A(n2704), .B(n11069), .C(n2680), .D(n6542), .Q(n8131) );
  OAI222 U1694 ( .A(n3040), .B(n11067), .C(n3016), .D(n6548), .Q(n8138) );
  OAI222 U1695 ( .A(n2992), .B(n11065), .C(n2968), .D(n6550), .Q(n8137) );
  OAI222 U1696 ( .A(n2944), .B(n11063), .C(n2920), .D(n6552), .Q(n8136) );
  OAI222 U1697 ( .A(n2896), .B(n11061), .C(n2872), .D(n6554), .Q(n8135) );
  OAI222 U1700 ( .A(n1696), .B(n11059), .C(n1672), .D(n6564), .Q(n8146) );
  OAI222 U1701 ( .A(n1648), .B(n11057), .C(n1624), .D(n6566), .Q(n8145) );
  OAI222 U1702 ( .A(n1600), .B(n11055), .C(n1576), .D(n6568), .Q(n8144) );
  OAI222 U1703 ( .A(n1552), .B(n11053), .C(n1528), .D(n6570), .Q(n8143) );
  OAI222 U1705 ( .A(n1888), .B(n11051), .C(n1864), .D(n6576), .Q(n8150) );
  OAI222 U1706 ( .A(n1840), .B(n11049), .C(n1816), .D(n6578), .Q(n8149) );
  OAI222 U1707 ( .A(n1792), .B(n11047), .C(n1768), .D(n6580), .Q(n8148) );
  OAI222 U1708 ( .A(n1744), .B(n11045), .C(n1720), .D(n6582), .Q(n8147) );
  OAI222 U1710 ( .A(n2080), .B(n11043), .C(n2056), .D(n6588), .Q(n8154) );
  OAI222 U1711 ( .A(n2032), .B(n11041), .C(n2008), .D(n6590), .Q(n8153) );
  OAI222 U1712 ( .A(n1984), .B(n11039), .C(n1960), .D(n6592), .Q(n8152) );
  OAI222 U1713 ( .A(n1936), .B(n11037), .C(n1912), .D(n6594), .Q(n8151) );
  OAI222 U1715 ( .A(n2272), .B(n11035), .C(n2248), .D(n6600), .Q(n8158) );
  OAI222 U1716 ( .A(n2224), .B(n11033), .C(n2200), .D(n6602), .Q(n8157) );
  OAI222 U1717 ( .A(n2176), .B(n11031), .C(n2152), .D(n6604), .Q(n8156) );
  OAI222 U1718 ( .A(n2128), .B(n11029), .C(n2104), .D(n6606), .Q(n8155) );
  OAI222 U1721 ( .A(n928), .B(n11027), .C(n904), .D(n6616), .Q(n8166) );
  OAI222 U1722 ( .A(n880), .B(n11025), .C(n856), .D(n6618), .Q(n8165) );
  OAI222 U1723 ( .A(n832), .B(n11023), .C(n808), .D(n6620), .Q(n8164) );
  OAI222 U1724 ( .A(n784), .B(n11021), .C(n760), .D(n6622), .Q(n8163) );
  OAI222 U1726 ( .A(n1120), .B(n11019), .C(n1096), .D(n6628), .Q(n8170) );
  OAI222 U1727 ( .A(n1072), .B(n11017), .C(n1048), .D(n6630), .Q(n8169) );
  OAI222 U1728 ( .A(n1024), .B(n11015), .C(n1000), .D(n6632), .Q(n8168) );
  OAI222 U1729 ( .A(n976), .B(n11013), .C(n952), .D(n6634), .Q(n8167) );
  OAI222 U1731 ( .A(n1312), .B(n11011), .C(n1288), .D(n6640), .Q(n8174) );
  OAI222 U1732 ( .A(n1264), .B(n11009), .C(n1240), .D(n6642), .Q(n8173) );
  OAI222 U1733 ( .A(n1216), .B(n11007), .C(n1192), .D(n6644), .Q(n8172) );
  OAI222 U1734 ( .A(n1168), .B(n11005), .C(n1144), .D(n6646), .Q(n8171) );
  OAI222 U1736 ( .A(n1504), .B(n11003), .C(n1480), .D(n6652), .Q(n8178) );
  OAI222 U1737 ( .A(n1456), .B(n11001), .C(n1432), .D(n6654), .Q(n8177) );
  OAI222 U1738 ( .A(n1408), .B(n10999), .C(n1384), .D(n6656), .Q(n8176) );
  OAI222 U1739 ( .A(n1360), .B(n10997), .C(n1336), .D(n6658), .Q(n8175) );
  OAI222 U1742 ( .A(n160), .B(n10995), .C(n136), .D(n6668), .Q(n8186) );
  OAI222 U1743 ( .A(n112), .B(n10993), .C(n88), .D(n6670), .Q(n8185) );
  OAI222 U1744 ( .A(n64), .B(n10991), .C(n40), .D(n6672), .Q(n8184) );
  OAI222 U1745 ( .A(n16), .B(n10989), .C(n6136), .D(n6674), .Q(n8183) );
  OAI222 U1747 ( .A(n352), .B(n10987), .C(n328), .D(n6680), .Q(n8190) );
  OAI222 U1748 ( .A(n304), .B(n10985), .C(n280), .D(n6682), .Q(n8189) );
  OAI222 U1749 ( .A(n256), .B(n10983), .C(n232), .D(n6684), .Q(n8188) );
  OAI222 U1750 ( .A(n208), .B(n10981), .C(n184), .D(n6686), .Q(n8187) );
  OAI222 U1752 ( .A(n544), .B(n10979), .C(n520), .D(n6692), .Q(n8194) );
  OAI222 U1753 ( .A(n496), .B(n10977), .C(n472), .D(n6694), .Q(n8193) );
  OAI222 U1754 ( .A(n448), .B(n10975), .C(n424), .D(n6696), .Q(n8192) );
  OAI222 U1755 ( .A(n400), .B(n10973), .C(n376), .D(n6698), .Q(n8191) );
  OAI222 U1757 ( .A(n736), .B(n10971), .C(n712), .D(n6704), .Q(n8198) );
  OAI222 U1758 ( .A(n688), .B(n10969), .C(n664), .D(n6706), .Q(n8197) );
  OAI222 U1759 ( .A(n640), .B(n10967), .C(n616), .D(n6708), .Q(n8196) );
  OAI222 U1760 ( .A(n592), .B(n10965), .C(n568), .D(n6710), .Q(n8195) );
  OAI222 U1764 ( .A(n5536), .B(n10963), .C(n5512), .D(n6724), .Q(n8210) );
  OAI222 U1765 ( .A(n5488), .B(n10961), .C(n5464), .D(n6726), .Q(n8209) );
  OAI222 U1766 ( .A(n5440), .B(n10959), .C(n5416), .D(n6728), .Q(n8208) );
  OAI222 U1767 ( .A(n5392), .B(n10957), .C(n5368), .D(n6730), .Q(n8207) );
  OAI222 U1769 ( .A(n5728), .B(n10955), .C(n5704), .D(n6736), .Q(n8214) );
  OAI222 U1770 ( .A(n5680), .B(n10953), .C(n5656), .D(n6738), .Q(n8213) );
  OAI222 U1771 ( .A(n5632), .B(n10951), .C(n5608), .D(n6740), .Q(n8212) );
  OAI222 U1772 ( .A(n5584), .B(n10949), .C(n5560), .D(n6742), .Q(n8211) );
  OAI222 U1774 ( .A(n5920), .B(n10947), .C(n5896), .D(n6748), .Q(n8218) );
  OAI222 U1775 ( .A(n5872), .B(n10945), .C(n5848), .D(n6750), .Q(n8217) );
  OAI222 U1776 ( .A(n5824), .B(n10943), .C(n5800), .D(n6752), .Q(n8216) );
  OAI222 U1777 ( .A(n5776), .B(n10941), .C(n5752), .D(n6754), .Q(n8215) );
  OAI222 U1779 ( .A(n6112), .B(n10939), .C(n6088), .D(n6760), .Q(n8222) );
  OAI222 U1780 ( .A(n6064), .B(n10937), .C(n6040), .D(n6762), .Q(n8221) );
  OAI222 U1781 ( .A(n6016), .B(n10935), .C(n5992), .D(n6764), .Q(n8220) );
  OAI222 U1782 ( .A(n5968), .B(n10933), .C(n5944), .D(n6766), .Q(n8219) );
  OAI222 U1785 ( .A(n4768), .B(n10931), .C(n4744), .D(n6776), .Q(n8230) );
  OAI222 U1786 ( .A(n4720), .B(n10929), .C(n4696), .D(n6778), .Q(n8229) );
  OAI222 U1787 ( .A(n4672), .B(n10927), .C(n4648), .D(n6780), .Q(n8228) );
  OAI222 U1788 ( .A(n4624), .B(n10925), .C(n4600), .D(n6782), .Q(n8227) );
  OAI222 U1790 ( .A(n4960), .B(n10923), .C(n4936), .D(n6788), .Q(n8234) );
  OAI222 U1791 ( .A(n4912), .B(n10921), .C(n4888), .D(n6790), .Q(n8233) );
  OAI222 U1792 ( .A(n4864), .B(n10919), .C(n4840), .D(n6792), .Q(n8232) );
  OAI222 U1793 ( .A(n4816), .B(n10917), .C(n4792), .D(n6794), .Q(n8231) );
  OAI222 U1795 ( .A(n5152), .B(n10915), .C(n5128), .D(n6800), .Q(n8238) );
  OAI222 U1796 ( .A(n5104), .B(n10913), .C(n5080), .D(n6802), .Q(n8237) );
  OAI222 U1797 ( .A(n5056), .B(n10911), .C(n5032), .D(n6804), .Q(n8236) );
  OAI222 U1798 ( .A(n5008), .B(n10909), .C(n4984), .D(n6806), .Q(n8235) );
  OAI222 U1800 ( .A(n5344), .B(n10907), .C(n5320), .D(n6812), .Q(n8242) );
  OAI222 U1801 ( .A(n5296), .B(n10905), .C(n5272), .D(n6814), .Q(n8241) );
  OAI222 U1802 ( .A(n5248), .B(n10903), .C(n5224), .D(n6816), .Q(n8240) );
  OAI222 U1803 ( .A(n5200), .B(n10901), .C(n5176), .D(n6818), .Q(n8239) );
  OAI222 U1806 ( .A(n4000), .B(n10899), .C(n3976), .D(n6828), .Q(n8250) );
  OAI222 U1807 ( .A(n3952), .B(n10897), .C(n3928), .D(n6830), .Q(n8249) );
  OAI222 U1808 ( .A(n3904), .B(n10895), .C(n3880), .D(n6832), .Q(n8248) );
  OAI222 U1809 ( .A(n3856), .B(n10893), .C(n3832), .D(n6834), .Q(n8247) );
  OAI222 U1811 ( .A(n4192), .B(n10891), .C(n4168), .D(n6840), .Q(n8254) );
  OAI222 U1812 ( .A(n4144), .B(n10889), .C(n4120), .D(n6842), .Q(n8253) );
  OAI222 U1813 ( .A(n4096), .B(n10887), .C(n4072), .D(n6844), .Q(n8252) );
  OAI222 U1814 ( .A(n4048), .B(n10885), .C(n4024), .D(n6846), .Q(n8251) );
  OAI222 U1816 ( .A(n4384), .B(n10883), .C(n4360), .D(n6852), .Q(n8258) );
  OAI222 U1817 ( .A(n4336), .B(n10881), .C(n4312), .D(n6854), .Q(n8257) );
  OAI222 U1818 ( .A(n4288), .B(n6191), .C(n4264), .D(n6856), .Q(n8256) );
  OAI222 U1819 ( .A(n4240), .B(n6189), .C(n4216), .D(n6858), .Q(n8255) );
  OAI222 U1821 ( .A(n4576), .B(n6187), .C(n4552), .D(n6864), .Q(n8262) );
  OAI222 U1822 ( .A(n4528), .B(n6185), .C(n4504), .D(n6866), .Q(n8261) );
  OAI222 U1823 ( .A(n4480), .B(n6183), .C(n4456), .D(n6868), .Q(n8260) );
  OAI222 U1824 ( .A(n4432), .B(n6181), .C(n4408), .D(n6870), .Q(n8259) );
  OAI222 U1827 ( .A(n3232), .B(n6179), .C(n3208), .D(n6880), .Q(n8270) );
  OAI222 U1828 ( .A(n3184), .B(n6177), .C(n3160), .D(n6882), .Q(n8269) );
  OAI222 U1829 ( .A(n3136), .B(n6175), .C(n3112), .D(n6884), .Q(n8268) );
  OAI222 U1830 ( .A(n3088), .B(n6173), .C(n3064), .D(n6886), .Q(n8267) );
  OAI222 U1832 ( .A(n3424), .B(n6171), .C(n3400), .D(n6892), .Q(n8274) );
  OAI222 U1833 ( .A(n3376), .B(n6169), .C(n3352), .D(n6894), .Q(n8273) );
  OAI222 U1834 ( .A(n3328), .B(n6167), .C(n3304), .D(n6896), .Q(n8272) );
  OAI222 U1835 ( .A(n3280), .B(n6165), .C(n3256), .D(n6898), .Q(n8271) );
  OAI222 U1837 ( .A(n3616), .B(n6163), .C(n3592), .D(n6904), .Q(n8278) );
  OAI222 U1838 ( .A(n3568), .B(n6161), .C(n3544), .D(n6906), .Q(n8277) );
  OAI222 U1839 ( .A(n3520), .B(n6159), .C(n3496), .D(n6908), .Q(n8276) );
  OAI222 U1840 ( .A(n3472), .B(n6157), .C(n3448), .D(n6910), .Q(n8275) );
  OAI222 U1842 ( .A(n3808), .B(n6155), .C(n3784), .D(n6916), .Q(n8282) );
  OAI222 U1843 ( .A(n3760), .B(n6153), .C(n3736), .D(n6918), .Q(n8281) );
  OAI222 U1844 ( .A(n3712), .B(n6151), .C(n3688), .D(n6920), .Q(n8280) );
  OAI222 U1845 ( .A(n3664), .B(n6149), .C(n3640), .D(n6922), .Q(n8279) );
  OAI222 U1850 ( .A(n2463), .B(n11091), .C(n2439), .D(n11297), .Q(n8296) );
  OAI222 U1851 ( .A(n2415), .B(n11089), .C(n2391), .D(n11296), .Q(n8295) );
  OAI222 U1852 ( .A(n2367), .B(n11087), .C(n2343), .D(n11295), .Q(n8294) );
  OAI222 U1853 ( .A(n2319), .B(n11085), .C(n2295), .D(n11294), .Q(n8293) );
  OAI222 U1855 ( .A(n2655), .B(n11083), .C(n2631), .D(n11293), .Q(n8300) );
  OAI222 U1856 ( .A(n2607), .B(n11081), .C(n2583), .D(n11292), .Q(n8299) );
  OAI222 U1857 ( .A(n2559), .B(n11079), .C(n2535), .D(n11291), .Q(n8298) );
  OAI222 U1858 ( .A(n2511), .B(n11077), .C(n2487), .D(n11290), .Q(n8297) );
  OAI222 U1860 ( .A(n2847), .B(n11075), .C(n2823), .D(n11289), .Q(n8304) );
  OAI222 U1861 ( .A(n2799), .B(n11073), .C(n2775), .D(n11288), .Q(n8303) );
  OAI222 U1862 ( .A(n2751), .B(n11071), .C(n2727), .D(n11287), .Q(n8302) );
  OAI222 U1863 ( .A(n2703), .B(n11069), .C(n2679), .D(n11286), .Q(n8301) );
  OAI222 U1865 ( .A(n3039), .B(n11067), .C(n3015), .D(n11285), .Q(n8308) );
  OAI222 U1866 ( .A(n2991), .B(n11065), .C(n2967), .D(n11284), .Q(n8307) );
  OAI222 U1867 ( .A(n2943), .B(n11063), .C(n2919), .D(n11283), .Q(n8306) );
  OAI222 U1868 ( .A(n2895), .B(n11061), .C(n2871), .D(n11282), .Q(n8305) );
  OAI222 U1871 ( .A(n1695), .B(n11059), .C(n1671), .D(n11281), .Q(n8316) );
  OAI222 U1872 ( .A(n1647), .B(n11057), .C(n1623), .D(n11280), .Q(n8315) );
  OAI222 U1873 ( .A(n1599), .B(n11055), .C(n1575), .D(n11279), .Q(n8314) );
  OAI222 U1874 ( .A(n1551), .B(n11053), .C(n1527), .D(n11278), .Q(n8313) );
  OAI222 U1876 ( .A(n1887), .B(n11051), .C(n1863), .D(n11277), .Q(n8320) );
  OAI222 U1877 ( .A(n1839), .B(n11049), .C(n1815), .D(n11276), .Q(n8319) );
  OAI222 U1878 ( .A(n1791), .B(n11047), .C(n1767), .D(n11275), .Q(n8318) );
  OAI222 U1879 ( .A(n1743), .B(n11045), .C(n1719), .D(n11274), .Q(n8317) );
  OAI222 U1881 ( .A(n2079), .B(n11043), .C(n2055), .D(n11273), .Q(n8324) );
  OAI222 U1882 ( .A(n2031), .B(n11041), .C(n2007), .D(n11272), .Q(n8323) );
  OAI222 U1883 ( .A(n1983), .B(n11039), .C(n1959), .D(n11271), .Q(n8322) );
  OAI222 U1884 ( .A(n1935), .B(n11037), .C(n1911), .D(n11270), .Q(n8321) );
  OAI222 U1886 ( .A(n2271), .B(n11035), .C(n2247), .D(n11269), .Q(n8328) );
  OAI222 U1887 ( .A(n2223), .B(n11033), .C(n2199), .D(n11268), .Q(n8327) );
  OAI222 U1888 ( .A(n2175), .B(n11031), .C(n2151), .D(n11267), .Q(n8326) );
  OAI222 U1889 ( .A(n2127), .B(n11029), .C(n2103), .D(n11266), .Q(n8325) );
  OAI222 U1892 ( .A(n927), .B(n11027), .C(n903), .D(n11265), .Q(n8336) );
  OAI222 U1893 ( .A(n879), .B(n11025), .C(n855), .D(n11264), .Q(n8335) );
  OAI222 U1894 ( .A(n831), .B(n11023), .C(n807), .D(n11263), .Q(n8334) );
  OAI222 U1895 ( .A(n783), .B(n11021), .C(n759), .D(n11262), .Q(n8333) );
  OAI222 U1897 ( .A(n1119), .B(n11019), .C(n1095), .D(n11261), .Q(n8340) );
  OAI222 U1898 ( .A(n1071), .B(n11017), .C(n1047), .D(n11260), .Q(n8339) );
  OAI222 U1899 ( .A(n1023), .B(n11015), .C(n999), .D(n11259), .Q(n8338) );
  OAI222 U1900 ( .A(n975), .B(n11013), .C(n951), .D(n11258), .Q(n8337) );
  OAI222 U1902 ( .A(n1311), .B(n11011), .C(n1287), .D(n11257), .Q(n8344) );
  OAI222 U1903 ( .A(n1263), .B(n11009), .C(n1239), .D(n11256), .Q(n8343) );
  OAI222 U1904 ( .A(n1215), .B(n11007), .C(n1191), .D(n11255), .Q(n8342) );
  OAI222 U1905 ( .A(n1167), .B(n11005), .C(n1143), .D(n11254), .Q(n8341) );
  OAI222 U1907 ( .A(n1503), .B(n11003), .C(n1479), .D(n11253), .Q(n8348) );
  OAI222 U1908 ( .A(n1455), .B(n11001), .C(n1431), .D(n11252), .Q(n8347) );
  OAI222 U1909 ( .A(n1407), .B(n10999), .C(n1383), .D(n11251), .Q(n8346) );
  OAI222 U1910 ( .A(n1359), .B(n10997), .C(n1335), .D(n11250), .Q(n8345) );
  OAI222 U1913 ( .A(n159), .B(n10995), .C(n135), .D(n11249), .Q(n8356) );
  OAI222 U1914 ( .A(n111), .B(n10993), .C(n87), .D(n11248), .Q(n8355) );
  OAI222 U1915 ( .A(n63), .B(n10991), .C(n39), .D(n11247), .Q(n8354) );
  OAI222 U1916 ( .A(n15), .B(n10989), .C(n6135), .D(n11246), .Q(n8353) );
  OAI222 U1918 ( .A(n351), .B(n10987), .C(n327), .D(n11245), .Q(n8360) );
  OAI222 U1919 ( .A(n303), .B(n10985), .C(n279), .D(n11244), .Q(n8359) );
  OAI222 U1920 ( .A(n255), .B(n10983), .C(n231), .D(n11243), .Q(n8358) );
  OAI222 U1921 ( .A(n207), .B(n10981), .C(n183), .D(n11242), .Q(n8357) );
  OAI222 U1923 ( .A(n543), .B(n10979), .C(n519), .D(n11241), .Q(n8364) );
  OAI222 U1924 ( .A(n495), .B(n10977), .C(n471), .D(n11240), .Q(n8363) );
  OAI222 U1925 ( .A(n447), .B(n10975), .C(n423), .D(n11239), .Q(n8362) );
  OAI222 U1926 ( .A(n399), .B(n10973), .C(n375), .D(n11238), .Q(n8361) );
  OAI222 U1928 ( .A(n735), .B(n10971), .C(n711), .D(n11237), .Q(n8368) );
  OAI222 U1929 ( .A(n687), .B(n10969), .C(n663), .D(n11236), .Q(n8367) );
  OAI222 U1930 ( .A(n639), .B(n10967), .C(n615), .D(n11235), .Q(n8366) );
  OAI222 U1931 ( .A(n591), .B(n10965), .C(n567), .D(n11234), .Q(n8365) );
  OAI222 U1935 ( .A(n5535), .B(n10963), .C(n5511), .D(n11233), .Q(n8380) );
  OAI222 U1936 ( .A(n5487), .B(n10961), .C(n5463), .D(n11232), .Q(n8379) );
  OAI222 U1937 ( .A(n5439), .B(n10959), .C(n5415), .D(n11231), .Q(n8378) );
  OAI222 U1938 ( .A(n5391), .B(n10957), .C(n5367), .D(n11230), .Q(n8377) );
  OAI222 U1940 ( .A(n5727), .B(n10955), .C(n5703), .D(n11229), .Q(n8384) );
  OAI222 U1941 ( .A(n5679), .B(n10953), .C(n5655), .D(n11228), .Q(n8383) );
  OAI222 U1942 ( .A(n5631), .B(n10951), .C(n5607), .D(n11227), .Q(n8382) );
  OAI222 U1943 ( .A(n5583), .B(n10949), .C(n5559), .D(n11226), .Q(n8381) );
  OAI222 U1945 ( .A(n5919), .B(n10947), .C(n5895), .D(n11225), .Q(n8388) );
  OAI222 U1946 ( .A(n5871), .B(n10945), .C(n5847), .D(n11224), .Q(n8387) );
  OAI222 U1947 ( .A(n5823), .B(n10943), .C(n5799), .D(n11223), .Q(n8386) );
  OAI222 U1948 ( .A(n5775), .B(n10941), .C(n5751), .D(n11222), .Q(n8385) );
  OAI222 U1950 ( .A(n6111), .B(n10939), .C(n6087), .D(n11221), .Q(n8392) );
  OAI222 U1951 ( .A(n6063), .B(n10937), .C(n6039), .D(n11220), .Q(n8391) );
  OAI222 U1952 ( .A(n6015), .B(n10935), .C(n5991), .D(n11219), .Q(n8390) );
  OAI222 U1953 ( .A(n5967), .B(n10933), .C(n5943), .D(n11218), .Q(n8389) );
  OAI222 U1956 ( .A(n4767), .B(n10931), .C(n4743), .D(n11217), .Q(n8400) );
  OAI222 U1957 ( .A(n4719), .B(n10929), .C(n4695), .D(n11216), .Q(n8399) );
  OAI222 U1958 ( .A(n4671), .B(n10927), .C(n4647), .D(n11215), .Q(n8398) );
  OAI222 U1959 ( .A(n4623), .B(n10925), .C(n4599), .D(n11214), .Q(n8397) );
  OAI222 U1961 ( .A(n4959), .B(n10923), .C(n4935), .D(n11213), .Q(n8404) );
  OAI222 U1962 ( .A(n4911), .B(n10921), .C(n4887), .D(n11212), .Q(n8403) );
  OAI222 U1963 ( .A(n4863), .B(n10919), .C(n4839), .D(n11211), .Q(n8402) );
  OAI222 U1964 ( .A(n4815), .B(n10917), .C(n4791), .D(n11210), .Q(n8401) );
  OAI222 U1966 ( .A(n5151), .B(n10915), .C(n5127), .D(n11209), .Q(n8408) );
  OAI222 U1967 ( .A(n5103), .B(n10913), .C(n5079), .D(n11208), .Q(n8407) );
  OAI222 U1968 ( .A(n5055), .B(n10911), .C(n5031), .D(n11207), .Q(n8406) );
  OAI222 U1969 ( .A(n5007), .B(n10909), .C(n4983), .D(n11206), .Q(n8405) );
  OAI222 U1971 ( .A(n5343), .B(n10907), .C(n5319), .D(n11205), .Q(n8412) );
  OAI222 U1972 ( .A(n5295), .B(n10905), .C(n5271), .D(n11204), .Q(n8411) );
  OAI222 U1973 ( .A(n5247), .B(n10903), .C(n5223), .D(n11203), .Q(n8410) );
  OAI222 U1974 ( .A(n5199), .B(n10901), .C(n5175), .D(n11202), .Q(n8409) );
  OAI222 U1977 ( .A(n3999), .B(n10899), .C(n3975), .D(n11201), .Q(n8420) );
  OAI222 U1978 ( .A(n3951), .B(n10897), .C(n3927), .D(n11200), .Q(n8419) );
  OAI222 U1979 ( .A(n3903), .B(n10895), .C(n3879), .D(n11199), .Q(n8418) );
  OAI222 U1980 ( .A(n3855), .B(n10893), .C(n3831), .D(n11198), .Q(n8417) );
  OAI222 U1982 ( .A(n4191), .B(n10891), .C(n4167), .D(n11197), .Q(n8424) );
  OAI222 U1983 ( .A(n4143), .B(n10889), .C(n4119), .D(n11196), .Q(n8423) );
  OAI222 U1984 ( .A(n4095), .B(n10887), .C(n4071), .D(n11195), .Q(n8422) );
  OAI222 U1985 ( .A(n4047), .B(n10885), .C(n4023), .D(n11194), .Q(n8421) );
  OAI222 U1987 ( .A(n4383), .B(n10883), .C(n4359), .D(n11193), .Q(n8428) );
  OAI222 U1988 ( .A(n4335), .B(n10881), .C(n4311), .D(n11192), .Q(n8427) );
  OAI222 U1989 ( .A(n4287), .B(n6191), .C(n4263), .D(n11191), .Q(n8426) );
  OAI222 U1990 ( .A(n4239), .B(n6189), .C(n4215), .D(n11190), .Q(n8425) );
  OAI222 U1992 ( .A(n4575), .B(n6187), .C(n4551), .D(n11189), .Q(n8432) );
  OAI222 U1993 ( .A(n4527), .B(n6185), .C(n4503), .D(n11188), .Q(n8431) );
  OAI222 U1994 ( .A(n4479), .B(n6183), .C(n4455), .D(n11187), .Q(n8430) );
  OAI222 U1995 ( .A(n4431), .B(n6181), .C(n4407), .D(n11186), .Q(n8429) );
  OAI222 U1998 ( .A(n3231), .B(n6179), .C(n3207), .D(n11185), .Q(n8440) );
  OAI222 U1999 ( .A(n3183), .B(n6177), .C(n3159), .D(n11184), .Q(n8439) );
  OAI222 U2000 ( .A(n3135), .B(n6175), .C(n3111), .D(n11183), .Q(n8438) );
  OAI222 U2001 ( .A(n3087), .B(n6173), .C(n3063), .D(n11182), .Q(n8437) );
  OAI222 U2003 ( .A(n3423), .B(n6171), .C(n3399), .D(n11181), .Q(n8444) );
  OAI222 U2004 ( .A(n3375), .B(n6169), .C(n3351), .D(n11180), .Q(n8443) );
  OAI222 U2005 ( .A(n3327), .B(n6167), .C(n3303), .D(n11179), .Q(n8442) );
  OAI222 U2006 ( .A(n3279), .B(n6165), .C(n3255), .D(n11178), .Q(n8441) );
  OAI222 U2008 ( .A(n3615), .B(n6163), .C(n3591), .D(n11177), .Q(n8448) );
  OAI222 U2009 ( .A(n3567), .B(n6161), .C(n3543), .D(n11176), .Q(n8447) );
  OAI222 U2010 ( .A(n3519), .B(n6159), .C(n3495), .D(n11175), .Q(n8446) );
  OAI222 U2011 ( .A(n3471), .B(n6157), .C(n3447), .D(n11174), .Q(n8445) );
  OAI222 U2013 ( .A(n3807), .B(n6155), .C(n3783), .D(n11173), .Q(n8452) );
  OAI222 U2014 ( .A(n3759), .B(n6153), .C(n3735), .D(n11172), .Q(n8451) );
  OAI222 U2015 ( .A(n3711), .B(n6151), .C(n3687), .D(n11171), .Q(n8450) );
  OAI222 U2016 ( .A(n3663), .B(n6149), .C(n3639), .D(n11170), .Q(n8449) );
  OAI222 U2021 ( .A(n2462), .B(n11091), .C(n2438), .D(n11297), .Q(n8466) );
  OAI222 U2022 ( .A(n2414), .B(n11089), .C(n2390), .D(n11296), .Q(n8465) );
  OAI222 U2023 ( .A(n2366), .B(n11087), .C(n2342), .D(n11295), .Q(n8464) );
  OAI222 U2024 ( .A(n2318), .B(n11085), .C(n2294), .D(n11294), .Q(n8463) );
  OAI222 U2026 ( .A(n2654), .B(n11083), .C(n2630), .D(n11293), .Q(n8470) );
  OAI222 U2027 ( .A(n2606), .B(n11081), .C(n2582), .D(n11292), .Q(n8469) );
  OAI222 U2028 ( .A(n2558), .B(n11079), .C(n2534), .D(n11291), .Q(n8468) );
  OAI222 U2029 ( .A(n2510), .B(n11077), .C(n2486), .D(n11290), .Q(n8467) );
  OAI222 U2031 ( .A(n2846), .B(n11075), .C(n2822), .D(n11289), .Q(n8474) );
  OAI222 U2032 ( .A(n2798), .B(n11073), .C(n2774), .D(n11288), .Q(n8473) );
  OAI222 U2033 ( .A(n2750), .B(n11071), .C(n2726), .D(n11287), .Q(n8472) );
  OAI222 U2034 ( .A(n2702), .B(n11069), .C(n2678), .D(n11286), .Q(n8471) );
  OAI222 U2036 ( .A(n3038), .B(n11067), .C(n3014), .D(n11285), .Q(n8478) );
  OAI222 U2037 ( .A(n2990), .B(n11065), .C(n2966), .D(n11284), .Q(n8477) );
  OAI222 U2038 ( .A(n2942), .B(n11063), .C(n2918), .D(n11283), .Q(n8476) );
  OAI222 U2039 ( .A(n2894), .B(n11061), .C(n2870), .D(n11282), .Q(n8475) );
  OAI222 U2042 ( .A(n1694), .B(n11059), .C(n1670), .D(n11281), .Q(n8486) );
  OAI222 U2043 ( .A(n1646), .B(n11057), .C(n1622), .D(n11280), .Q(n8485) );
  OAI222 U2044 ( .A(n1598), .B(n11055), .C(n1574), .D(n11279), .Q(n8484) );
  OAI222 U2045 ( .A(n1550), .B(n11053), .C(n1526), .D(n11278), .Q(n8483) );
  OAI222 U2047 ( .A(n1886), .B(n11051), .C(n1862), .D(n11277), .Q(n8490) );
  OAI222 U2048 ( .A(n1838), .B(n11049), .C(n1814), .D(n11276), .Q(n8489) );
  OAI222 U2049 ( .A(n1790), .B(n11047), .C(n1766), .D(n11275), .Q(n8488) );
  OAI222 U2050 ( .A(n1742), .B(n11045), .C(n1718), .D(n11274), .Q(n8487) );
  OAI222 U2052 ( .A(n2078), .B(n11043), .C(n2054), .D(n11273), .Q(n8494) );
  OAI222 U2053 ( .A(n2030), .B(n11041), .C(n2006), .D(n11272), .Q(n8493) );
  OAI222 U2054 ( .A(n1982), .B(n11039), .C(n1958), .D(n11271), .Q(n8492) );
  OAI222 U2055 ( .A(n1934), .B(n11037), .C(n1910), .D(n11270), .Q(n8491) );
  OAI222 U2057 ( .A(n2270), .B(n11035), .C(n2246), .D(n11269), .Q(n8498) );
  OAI222 U2058 ( .A(n2222), .B(n11033), .C(n2198), .D(n11268), .Q(n8497) );
  OAI222 U2059 ( .A(n2174), .B(n11031), .C(n2150), .D(n11267), .Q(n8496) );
  OAI222 U2060 ( .A(n2126), .B(n11029), .C(n2102), .D(n11266), .Q(n8495) );
  OAI222 U2063 ( .A(n926), .B(n11027), .C(n902), .D(n11265), .Q(n8506) );
  OAI222 U2064 ( .A(n878), .B(n11025), .C(n854), .D(n11264), .Q(n8505) );
  OAI222 U2065 ( .A(n830), .B(n11023), .C(n806), .D(n11263), .Q(n8504) );
  OAI222 U2066 ( .A(n782), .B(n11021), .C(n758), .D(n11262), .Q(n8503) );
  OAI222 U2068 ( .A(n1118), .B(n11019), .C(n1094), .D(n11261), .Q(n8510) );
  OAI222 U2069 ( .A(n1070), .B(n11017), .C(n1046), .D(n11260), .Q(n8509) );
  OAI222 U2070 ( .A(n1022), .B(n11015), .C(n998), .D(n11259), .Q(n8508) );
  OAI222 U2071 ( .A(n974), .B(n11013), .C(n950), .D(n11258), .Q(n8507) );
  OAI222 U2073 ( .A(n1310), .B(n11011), .C(n1286), .D(n11257), .Q(n8514) );
  OAI222 U2074 ( .A(n1262), .B(n11009), .C(n1238), .D(n11256), .Q(n8513) );
  OAI222 U2075 ( .A(n1214), .B(n11007), .C(n1190), .D(n11255), .Q(n8512) );
  OAI222 U2076 ( .A(n1166), .B(n11005), .C(n1142), .D(n11254), .Q(n8511) );
  OAI222 U2078 ( .A(n1502), .B(n11003), .C(n1478), .D(n11253), .Q(n8518) );
  OAI222 U2079 ( .A(n1454), .B(n11001), .C(n1430), .D(n11252), .Q(n8517) );
  OAI222 U2080 ( .A(n1406), .B(n10999), .C(n1382), .D(n11251), .Q(n8516) );
  OAI222 U2081 ( .A(n1358), .B(n10997), .C(n1334), .D(n11250), .Q(n8515) );
  OAI222 U2084 ( .A(n158), .B(n10995), .C(n134), .D(n11249), .Q(n8526) );
  OAI222 U2085 ( .A(n110), .B(n10993), .C(n86), .D(n11248), .Q(n8525) );
  OAI222 U2086 ( .A(n62), .B(n10991), .C(n38), .D(n11247), .Q(n8524) );
  OAI222 U2087 ( .A(n14), .B(n10989), .C(n6134), .D(n11246), .Q(n8523) );
  OAI222 U2089 ( .A(n350), .B(n10987), .C(n326), .D(n11245), .Q(n8530) );
  OAI222 U2090 ( .A(n302), .B(n10985), .C(n278), .D(n11244), .Q(n8529) );
  OAI222 U2091 ( .A(n254), .B(n10983), .C(n230), .D(n11243), .Q(n8528) );
  OAI222 U2092 ( .A(n206), .B(n10981), .C(n182), .D(n11242), .Q(n8527) );
  OAI222 U2094 ( .A(n542), .B(n10979), .C(n518), .D(n11241), .Q(n8534) );
  OAI222 U2095 ( .A(n494), .B(n10977), .C(n470), .D(n11240), .Q(n8533) );
  OAI222 U2096 ( .A(n446), .B(n10975), .C(n422), .D(n11239), .Q(n8532) );
  OAI222 U2097 ( .A(n398), .B(n10973), .C(n374), .D(n11238), .Q(n8531) );
  OAI222 U2099 ( .A(n734), .B(n10971), .C(n710), .D(n11237), .Q(n8538) );
  OAI222 U2100 ( .A(n686), .B(n10969), .C(n662), .D(n11236), .Q(n8537) );
  OAI222 U2101 ( .A(n638), .B(n10967), .C(n614), .D(n11235), .Q(n8536) );
  OAI222 U2102 ( .A(n590), .B(n10965), .C(n566), .D(n11234), .Q(n8535) );
  OAI222 U2106 ( .A(n5534), .B(n10963), .C(n5510), .D(n11233), .Q(n8550) );
  OAI222 U2107 ( .A(n5486), .B(n10961), .C(n5462), .D(n11232), .Q(n8549) );
  OAI222 U2108 ( .A(n5438), .B(n10959), .C(n5414), .D(n11231), .Q(n8548) );
  OAI222 U2109 ( .A(n5390), .B(n10957), .C(n5366), .D(n11230), .Q(n8547) );
  OAI222 U2111 ( .A(n5726), .B(n10955), .C(n5702), .D(n11229), .Q(n8554) );
  OAI222 U2112 ( .A(n5678), .B(n10953), .C(n5654), .D(n11228), .Q(n8553) );
  OAI222 U2113 ( .A(n5630), .B(n10951), .C(n5606), .D(n11227), .Q(n8552) );
  OAI222 U2114 ( .A(n5582), .B(n10949), .C(n5558), .D(n11226), .Q(n8551) );
  OAI222 U2116 ( .A(n5918), .B(n10947), .C(n5894), .D(n11225), .Q(n8558) );
  OAI222 U2117 ( .A(n5870), .B(n10945), .C(n5846), .D(n11224), .Q(n8557) );
  OAI222 U2118 ( .A(n5822), .B(n10943), .C(n5798), .D(n11223), .Q(n8556) );
  OAI222 U2119 ( .A(n5774), .B(n10941), .C(n5750), .D(n11222), .Q(n8555) );
  OAI222 U2121 ( .A(n6110), .B(n10939), .C(n6086), .D(n11221), .Q(n8562) );
  OAI222 U2122 ( .A(n6062), .B(n10937), .C(n6038), .D(n11220), .Q(n8561) );
  OAI222 U2123 ( .A(n6014), .B(n10935), .C(n5990), .D(n11219), .Q(n8560) );
  OAI222 U2124 ( .A(n5966), .B(n10933), .C(n5942), .D(n11218), .Q(n8559) );
  OAI222 U2127 ( .A(n4766), .B(n10931), .C(n4742), .D(n11217), .Q(n8570) );
  OAI222 U2128 ( .A(n4718), .B(n10929), .C(n4694), .D(n11216), .Q(n8569) );
  OAI222 U2129 ( .A(n4670), .B(n10927), .C(n4646), .D(n11215), .Q(n8568) );
  OAI222 U2130 ( .A(n4622), .B(n10925), .C(n4598), .D(n11214), .Q(n8567) );
  OAI222 U2132 ( .A(n4958), .B(n10923), .C(n4934), .D(n11213), .Q(n8574) );
  OAI222 U2133 ( .A(n4910), .B(n10921), .C(n4886), .D(n11212), .Q(n8573) );
  OAI222 U2134 ( .A(n4862), .B(n10919), .C(n4838), .D(n11211), .Q(n8572) );
  OAI222 U2135 ( .A(n4814), .B(n10917), .C(n4790), .D(n11210), .Q(n8571) );
  OAI222 U2137 ( .A(n5150), .B(n10915), .C(n5126), .D(n11209), .Q(n8578) );
  OAI222 U2138 ( .A(n5102), .B(n10913), .C(n5078), .D(n11208), .Q(n8577) );
  OAI222 U2139 ( .A(n5054), .B(n10911), .C(n5030), .D(n11207), .Q(n8576) );
  OAI222 U2140 ( .A(n5006), .B(n10909), .C(n4982), .D(n11206), .Q(n8575) );
  OAI222 U2142 ( .A(n5342), .B(n10907), .C(n5318), .D(n11205), .Q(n8582) );
  OAI222 U2143 ( .A(n5294), .B(n10905), .C(n5270), .D(n11204), .Q(n8581) );
  OAI222 U2144 ( .A(n5246), .B(n10903), .C(n5222), .D(n11203), .Q(n8580) );
  OAI222 U2145 ( .A(n5198), .B(n10901), .C(n5174), .D(n11202), .Q(n8579) );
  OAI222 U2148 ( .A(n3998), .B(n10899), .C(n3974), .D(n11201), .Q(n8590) );
  OAI222 U2149 ( .A(n3950), .B(n10897), .C(n3926), .D(n11200), .Q(n8589) );
  OAI222 U2150 ( .A(n3902), .B(n10895), .C(n3878), .D(n11199), .Q(n8588) );
  OAI222 U2151 ( .A(n3854), .B(n10893), .C(n3830), .D(n11198), .Q(n8587) );
  OAI222 U2153 ( .A(n4190), .B(n10891), .C(n4166), .D(n11197), .Q(n8594) );
  OAI222 U2154 ( .A(n4142), .B(n10889), .C(n4118), .D(n11196), .Q(n8593) );
  OAI222 U2155 ( .A(n4094), .B(n10887), .C(n4070), .D(n11195), .Q(n8592) );
  OAI222 U2156 ( .A(n4046), .B(n10885), .C(n4022), .D(n11194), .Q(n8591) );
  OAI222 U2158 ( .A(n4382), .B(n10883), .C(n4358), .D(n11193), .Q(n8598) );
  OAI222 U2159 ( .A(n4334), .B(n10881), .C(n4310), .D(n11192), .Q(n8597) );
  OAI222 U2160 ( .A(n4286), .B(n6191), .C(n4262), .D(n11191), .Q(n8596) );
  OAI222 U2161 ( .A(n4238), .B(n6189), .C(n4214), .D(n11190), .Q(n8595) );
  OAI222 U2163 ( .A(n4574), .B(n6187), .C(n4550), .D(n11189), .Q(n8602) );
  OAI222 U2164 ( .A(n4526), .B(n6185), .C(n4502), .D(n11188), .Q(n8601) );
  OAI222 U2165 ( .A(n4478), .B(n6183), .C(n4454), .D(n11187), .Q(n8600) );
  OAI222 U2166 ( .A(n4430), .B(n6181), .C(n4406), .D(n11186), .Q(n8599) );
  OAI222 U2169 ( .A(n3230), .B(n6179), .C(n3206), .D(n11185), .Q(n8610) );
  OAI222 U2170 ( .A(n3182), .B(n6177), .C(n3158), .D(n11184), .Q(n8609) );
  OAI222 U2171 ( .A(n3134), .B(n6175), .C(n3110), .D(n11183), .Q(n8608) );
  OAI222 U2172 ( .A(n3086), .B(n6173), .C(n3062), .D(n11182), .Q(n8607) );
  OAI222 U2174 ( .A(n3422), .B(n6171), .C(n3398), .D(n11181), .Q(n8614) );
  OAI222 U2175 ( .A(n3374), .B(n6169), .C(n3350), .D(n11180), .Q(n8613) );
  OAI222 U2176 ( .A(n3326), .B(n6167), .C(n3302), .D(n11179), .Q(n8612) );
  OAI222 U2177 ( .A(n3278), .B(n6165), .C(n3254), .D(n11178), .Q(n8611) );
  OAI222 U2179 ( .A(n3614), .B(n6163), .C(n3590), .D(n11177), .Q(n8618) );
  OAI222 U2180 ( .A(n3566), .B(n6161), .C(n3542), .D(n11176), .Q(n8617) );
  OAI222 U2181 ( .A(n3518), .B(n6159), .C(n3494), .D(n11175), .Q(n8616) );
  OAI222 U2182 ( .A(n3470), .B(n6157), .C(n3446), .D(n11174), .Q(n8615) );
  OAI222 U2184 ( .A(n3806), .B(n6155), .C(n3782), .D(n11173), .Q(n8622) );
  OAI222 U2185 ( .A(n3758), .B(n6153), .C(n3734), .D(n11172), .Q(n8621) );
  OAI222 U2186 ( .A(n3710), .B(n6151), .C(n3686), .D(n11171), .Q(n8620) );
  OAI222 U2187 ( .A(n3662), .B(n6149), .C(n3638), .D(n11170), .Q(n8619) );
  OAI222 U2192 ( .A(n2461), .B(n11091), .C(n2437), .D(n11297), .Q(n8636) );
  OAI222 U2193 ( .A(n2413), .B(n11089), .C(n2389), .D(n11296), .Q(n8635) );
  OAI222 U2194 ( .A(n2365), .B(n11087), .C(n2341), .D(n11295), .Q(n8634) );
  OAI222 U2195 ( .A(n2317), .B(n11085), .C(n2293), .D(n11294), .Q(n8633) );
  OAI222 U2197 ( .A(n2653), .B(n11083), .C(n2629), .D(n11293), .Q(n8640) );
  OAI222 U2198 ( .A(n2605), .B(n11081), .C(n2581), .D(n11292), .Q(n8639) );
  OAI222 U2199 ( .A(n2557), .B(n11079), .C(n2533), .D(n11291), .Q(n8638) );
  OAI222 U2200 ( .A(n2509), .B(n11077), .C(n2485), .D(n11290), .Q(n8637) );
  OAI222 U2202 ( .A(n2845), .B(n11075), .C(n2821), .D(n11289), .Q(n8644) );
  OAI222 U2203 ( .A(n2797), .B(n11073), .C(n2773), .D(n11288), .Q(n8643) );
  OAI222 U2204 ( .A(n2749), .B(n11071), .C(n2725), .D(n11287), .Q(n8642) );
  OAI222 U2205 ( .A(n2701), .B(n11069), .C(n2677), .D(n11286), .Q(n8641) );
  OAI222 U2207 ( .A(n3037), .B(n11067), .C(n3013), .D(n11285), .Q(n8648) );
  OAI222 U2208 ( .A(n2989), .B(n11065), .C(n2965), .D(n11284), .Q(n8647) );
  OAI222 U2209 ( .A(n2941), .B(n11063), .C(n2917), .D(n11283), .Q(n8646) );
  OAI222 U2210 ( .A(n2893), .B(n11061), .C(n2869), .D(n11282), .Q(n8645) );
  OAI222 U2213 ( .A(n1693), .B(n11059), .C(n1669), .D(n11281), .Q(n8656) );
  OAI222 U2214 ( .A(n1645), .B(n11057), .C(n1621), .D(n11280), .Q(n8655) );
  OAI222 U2215 ( .A(n1597), .B(n11055), .C(n1573), .D(n11279), .Q(n8654) );
  OAI222 U2216 ( .A(n1549), .B(n11053), .C(n1525), .D(n11278), .Q(n8653) );
  OAI222 U2218 ( .A(n1885), .B(n11051), .C(n1861), .D(n11277), .Q(n8660) );
  OAI222 U2219 ( .A(n1837), .B(n11049), .C(n1813), .D(n11276), .Q(n8659) );
  OAI222 U2220 ( .A(n1789), .B(n11047), .C(n1765), .D(n11275), .Q(n8658) );
  OAI222 U2221 ( .A(n1741), .B(n11045), .C(n1717), .D(n11274), .Q(n8657) );
  OAI222 U2223 ( .A(n2077), .B(n11043), .C(n2053), .D(n11273), .Q(n8664) );
  OAI222 U2224 ( .A(n2029), .B(n11041), .C(n2005), .D(n11272), .Q(n8663) );
  OAI222 U2225 ( .A(n1981), .B(n11039), .C(n1957), .D(n11271), .Q(n8662) );
  OAI222 U2226 ( .A(n1933), .B(n11037), .C(n1909), .D(n11270), .Q(n8661) );
  OAI222 U2228 ( .A(n2269), .B(n11035), .C(n2245), .D(n11269), .Q(n8668) );
  OAI222 U2229 ( .A(n2221), .B(n11033), .C(n2197), .D(n11268), .Q(n8667) );
  OAI222 U2230 ( .A(n2173), .B(n11031), .C(n2149), .D(n11267), .Q(n8666) );
  OAI222 U2231 ( .A(n2125), .B(n11029), .C(n2101), .D(n11266), .Q(n8665) );
  OAI222 U2234 ( .A(n925), .B(n11027), .C(n901), .D(n11265), .Q(n8676) );
  OAI222 U2235 ( .A(n877), .B(n11025), .C(n853), .D(n11264), .Q(n8675) );
  OAI222 U2236 ( .A(n829), .B(n11023), .C(n805), .D(n11263), .Q(n8674) );
  OAI222 U2237 ( .A(n781), .B(n11021), .C(n757), .D(n11262), .Q(n8673) );
  OAI222 U2239 ( .A(n1117), .B(n11019), .C(n1093), .D(n11261), .Q(n8680) );
  OAI222 U2240 ( .A(n1069), .B(n11017), .C(n1045), .D(n11260), .Q(n8679) );
  OAI222 U2241 ( .A(n1021), .B(n11015), .C(n997), .D(n11259), .Q(n8678) );
  OAI222 U2242 ( .A(n973), .B(n11013), .C(n949), .D(n11258), .Q(n8677) );
  OAI222 U2244 ( .A(n1309), .B(n11011), .C(n1285), .D(n11257), .Q(n8684) );
  OAI222 U2245 ( .A(n1261), .B(n11009), .C(n1237), .D(n11256), .Q(n8683) );
  OAI222 U2246 ( .A(n1213), .B(n11007), .C(n1189), .D(n11255), .Q(n8682) );
  OAI222 U2247 ( .A(n1165), .B(n11005), .C(n1141), .D(n11254), .Q(n8681) );
  OAI222 U2249 ( .A(n1501), .B(n11003), .C(n1477), .D(n11253), .Q(n8688) );
  OAI222 U2250 ( .A(n1453), .B(n11001), .C(n1429), .D(n11252), .Q(n8687) );
  OAI222 U2251 ( .A(n1405), .B(n10999), .C(n1381), .D(n11251), .Q(n8686) );
  OAI222 U2252 ( .A(n1357), .B(n10997), .C(n1333), .D(n11250), .Q(n8685) );
  OAI222 U2255 ( .A(n157), .B(n10995), .C(n133), .D(n11249), .Q(n8696) );
  OAI222 U2256 ( .A(n109), .B(n10993), .C(n85), .D(n11248), .Q(n8695) );
  OAI222 U2257 ( .A(n61), .B(n10991), .C(n37), .D(n11247), .Q(n8694) );
  OAI222 U2258 ( .A(n13), .B(n10989), .C(n6133), .D(n11246), .Q(n8693) );
  OAI222 U2260 ( .A(n349), .B(n10987), .C(n325), .D(n11245), .Q(n8700) );
  OAI222 U2261 ( .A(n301), .B(n10985), .C(n277), .D(n11244), .Q(n8699) );
  OAI222 U2262 ( .A(n253), .B(n10983), .C(n229), .D(n11243), .Q(n8698) );
  OAI222 U2263 ( .A(n205), .B(n10981), .C(n181), .D(n11242), .Q(n8697) );
  OAI222 U2265 ( .A(n541), .B(n10979), .C(n517), .D(n11241), .Q(n8704) );
  OAI222 U2266 ( .A(n493), .B(n10977), .C(n469), .D(n11240), .Q(n8703) );
  OAI222 U2267 ( .A(n445), .B(n10975), .C(n421), .D(n11239), .Q(n8702) );
  OAI222 U2268 ( .A(n397), .B(n10973), .C(n373), .D(n11238), .Q(n8701) );
  OAI222 U2270 ( .A(n733), .B(n10971), .C(n709), .D(n11237), .Q(n8708) );
  OAI222 U2271 ( .A(n685), .B(n10969), .C(n661), .D(n11236), .Q(n8707) );
  OAI222 U2272 ( .A(n637), .B(n10967), .C(n613), .D(n11235), .Q(n8706) );
  OAI222 U2273 ( .A(n589), .B(n10965), .C(n565), .D(n11234), .Q(n8705) );
  OAI222 U2277 ( .A(n5533), .B(n10963), .C(n5509), .D(n11233), .Q(n8720) );
  OAI222 U2278 ( .A(n5485), .B(n10961), .C(n5461), .D(n11232), .Q(n8719) );
  OAI222 U2279 ( .A(n5437), .B(n10959), .C(n5413), .D(n11231), .Q(n8718) );
  OAI222 U2280 ( .A(n5389), .B(n10957), .C(n5365), .D(n11230), .Q(n8717) );
  OAI222 U2282 ( .A(n5725), .B(n10955), .C(n5701), .D(n11229), .Q(n8724) );
  OAI222 U2283 ( .A(n5677), .B(n10953), .C(n5653), .D(n11228), .Q(n8723) );
  OAI222 U2284 ( .A(n5629), .B(n10951), .C(n5605), .D(n11227), .Q(n8722) );
  OAI222 U2285 ( .A(n5581), .B(n10949), .C(n5557), .D(n11226), .Q(n8721) );
  OAI222 U2287 ( .A(n5917), .B(n10947), .C(n5893), .D(n11225), .Q(n8728) );
  OAI222 U2288 ( .A(n5869), .B(n10945), .C(n5845), .D(n11224), .Q(n8727) );
  OAI222 U2289 ( .A(n5821), .B(n10943), .C(n5797), .D(n11223), .Q(n8726) );
  OAI222 U2290 ( .A(n5773), .B(n10941), .C(n5749), .D(n11222), .Q(n8725) );
  OAI222 U2292 ( .A(n6109), .B(n10939), .C(n6085), .D(n11221), .Q(n8732) );
  OAI222 U2293 ( .A(n6061), .B(n10937), .C(n6037), .D(n11220), .Q(n8731) );
  OAI222 U2294 ( .A(n6013), .B(n10935), .C(n5989), .D(n11219), .Q(n8730) );
  OAI222 U2295 ( .A(n5965), .B(n10933), .C(n5941), .D(n11218), .Q(n8729) );
  OAI222 U2298 ( .A(n4765), .B(n10931), .C(n4741), .D(n11217), .Q(n8740) );
  OAI222 U2299 ( .A(n4717), .B(n10929), .C(n4693), .D(n11216), .Q(n8739) );
  OAI222 U2300 ( .A(n4669), .B(n10927), .C(n4645), .D(n11215), .Q(n8738) );
  OAI222 U2301 ( .A(n4621), .B(n10925), .C(n4597), .D(n11214), .Q(n8737) );
  OAI222 U2303 ( .A(n4957), .B(n10923), .C(n4933), .D(n11213), .Q(n8744) );
  OAI222 U2304 ( .A(n4909), .B(n10921), .C(n4885), .D(n11212), .Q(n8743) );
  OAI222 U2305 ( .A(n4861), .B(n10919), .C(n4837), .D(n11211), .Q(n8742) );
  OAI222 U2306 ( .A(n4813), .B(n10917), .C(n4789), .D(n11210), .Q(n8741) );
  OAI222 U2308 ( .A(n5149), .B(n10915), .C(n5125), .D(n11209), .Q(n8748) );
  OAI222 U2309 ( .A(n5101), .B(n10913), .C(n5077), .D(n11208), .Q(n8747) );
  OAI222 U2310 ( .A(n5053), .B(n10911), .C(n5029), .D(n11207), .Q(n8746) );
  OAI222 U2311 ( .A(n5005), .B(n10909), .C(n4981), .D(n11206), .Q(n8745) );
  OAI222 U2313 ( .A(n5341), .B(n10907), .C(n5317), .D(n11205), .Q(n8752) );
  OAI222 U2314 ( .A(n5293), .B(n10905), .C(n5269), .D(n11204), .Q(n8751) );
  OAI222 U2315 ( .A(n5245), .B(n10903), .C(n5221), .D(n11203), .Q(n8750) );
  OAI222 U2316 ( .A(n5197), .B(n10901), .C(n5173), .D(n11202), .Q(n8749) );
  OAI222 U2319 ( .A(n3997), .B(n10899), .C(n3973), .D(n11201), .Q(n8760) );
  OAI222 U2320 ( .A(n3949), .B(n10897), .C(n3925), .D(n11200), .Q(n8759) );
  OAI222 U2321 ( .A(n3901), .B(n10895), .C(n3877), .D(n11199), .Q(n8758) );
  OAI222 U2322 ( .A(n3853), .B(n10893), .C(n3829), .D(n11198), .Q(n8757) );
  OAI222 U2324 ( .A(n4189), .B(n10891), .C(n4165), .D(n11197), .Q(n8764) );
  OAI222 U2325 ( .A(n4141), .B(n10889), .C(n4117), .D(n11196), .Q(n8763) );
  OAI222 U2326 ( .A(n4093), .B(n10887), .C(n4069), .D(n11195), .Q(n8762) );
  OAI222 U2327 ( .A(n4045), .B(n10885), .C(n4021), .D(n11194), .Q(n8761) );
  OAI222 U2329 ( .A(n4381), .B(n10883), .C(n4357), .D(n11193), .Q(n8768) );
  OAI222 U2330 ( .A(n4333), .B(n10881), .C(n4309), .D(n11192), .Q(n8767) );
  OAI222 U2331 ( .A(n4285), .B(n6191), .C(n4261), .D(n11191), .Q(n8766) );
  OAI222 U2332 ( .A(n4237), .B(n6189), .C(n4213), .D(n11190), .Q(n8765) );
  OAI222 U2334 ( .A(n4573), .B(n6187), .C(n4549), .D(n11189), .Q(n8772) );
  OAI222 U2335 ( .A(n4525), .B(n6185), .C(n4501), .D(n11188), .Q(n8771) );
  OAI222 U2336 ( .A(n4477), .B(n6183), .C(n4453), .D(n11187), .Q(n8770) );
  OAI222 U2337 ( .A(n4429), .B(n6181), .C(n4405), .D(n11186), .Q(n8769) );
  OAI222 U2340 ( .A(n3229), .B(n6179), .C(n3205), .D(n11185), .Q(n8780) );
  OAI222 U2341 ( .A(n3181), .B(n6177), .C(n3157), .D(n11184), .Q(n8779) );
  OAI222 U2342 ( .A(n3133), .B(n6175), .C(n3109), .D(n11183), .Q(n8778) );
  OAI222 U2343 ( .A(n3085), .B(n6173), .C(n3061), .D(n11182), .Q(n8777) );
  OAI222 U2345 ( .A(n3421), .B(n6171), .C(n3397), .D(n11181), .Q(n8784) );
  OAI222 U2346 ( .A(n3373), .B(n6169), .C(n3349), .D(n11180), .Q(n8783) );
  OAI222 U2347 ( .A(n3325), .B(n6167), .C(n3301), .D(n11179), .Q(n8782) );
  OAI222 U2348 ( .A(n3277), .B(n6165), .C(n3253), .D(n11178), .Q(n8781) );
  OAI222 U2350 ( .A(n3613), .B(n6163), .C(n3589), .D(n11177), .Q(n8788) );
  OAI222 U2351 ( .A(n3565), .B(n6161), .C(n3541), .D(n11176), .Q(n8787) );
  OAI222 U2352 ( .A(n3517), .B(n6159), .C(n3493), .D(n11175), .Q(n8786) );
  OAI222 U2353 ( .A(n3469), .B(n6157), .C(n3445), .D(n11174), .Q(n8785) );
  OAI222 U2355 ( .A(n3805), .B(n6155), .C(n3781), .D(n11173), .Q(n8792) );
  OAI222 U2356 ( .A(n3757), .B(n6153), .C(n3733), .D(n11172), .Q(n8791) );
  OAI222 U2357 ( .A(n3709), .B(n6151), .C(n3685), .D(n11171), .Q(n8790) );
  OAI222 U2358 ( .A(n3661), .B(n6149), .C(n3637), .D(n11170), .Q(n8789) );
  OAI222 U2363 ( .A(n2460), .B(n11090), .C(n2436), .D(n11297), .Q(n8806) );
  OAI222 U2364 ( .A(n2412), .B(n11088), .C(n2388), .D(n11296), .Q(n8805) );
  OAI222 U2365 ( .A(n2364), .B(n11086), .C(n2340), .D(n11295), .Q(n8804) );
  OAI222 U2366 ( .A(n2316), .B(n11084), .C(n2292), .D(n11294), .Q(n8803) );
  OAI222 U2368 ( .A(n2652), .B(n11082), .C(n2628), .D(n11293), .Q(n8810) );
  OAI222 U2369 ( .A(n2604), .B(n11080), .C(n2580), .D(n11292), .Q(n8809) );
  OAI222 U2370 ( .A(n2556), .B(n11078), .C(n2532), .D(n11291), .Q(n8808) );
  OAI222 U2371 ( .A(n2508), .B(n11076), .C(n2484), .D(n11290), .Q(n8807) );
  OAI222 U2373 ( .A(n2844), .B(n11074), .C(n2820), .D(n11289), .Q(n8814) );
  OAI222 U2374 ( .A(n2796), .B(n11072), .C(n2772), .D(n11288), .Q(n8813) );
  OAI222 U2375 ( .A(n2748), .B(n11070), .C(n2724), .D(n11287), .Q(n8812) );
  OAI222 U2376 ( .A(n2700), .B(n11068), .C(n2676), .D(n11286), .Q(n8811) );
  OAI222 U2378 ( .A(n3036), .B(n11066), .C(n3012), .D(n11285), .Q(n8818) );
  OAI222 U2379 ( .A(n2988), .B(n11064), .C(n2964), .D(n11284), .Q(n8817) );
  OAI222 U2380 ( .A(n2940), .B(n11062), .C(n2916), .D(n11283), .Q(n8816) );
  OAI222 U2381 ( .A(n2892), .B(n11060), .C(n2868), .D(n11282), .Q(n8815) );
  OAI222 U2384 ( .A(n1692), .B(n11058), .C(n1668), .D(n11281), .Q(n8826) );
  OAI222 U2385 ( .A(n1644), .B(n11056), .C(n1620), .D(n11280), .Q(n8825) );
  OAI222 U2386 ( .A(n1596), .B(n11054), .C(n1572), .D(n11279), .Q(n8824) );
  OAI222 U2387 ( .A(n1548), .B(n11052), .C(n1524), .D(n11278), .Q(n8823) );
  OAI222 U2389 ( .A(n1884), .B(n11050), .C(n1860), .D(n11277), .Q(n8830) );
  OAI222 U2390 ( .A(n1836), .B(n11048), .C(n1812), .D(n11276), .Q(n8829) );
  OAI222 U2391 ( .A(n1788), .B(n11046), .C(n1764), .D(n11275), .Q(n8828) );
  OAI222 U2392 ( .A(n1740), .B(n11044), .C(n1716), .D(n11274), .Q(n8827) );
  OAI222 U2394 ( .A(n2076), .B(n11042), .C(n2052), .D(n11273), .Q(n8834) );
  OAI222 U2395 ( .A(n2028), .B(n11040), .C(n2004), .D(n11272), .Q(n8833) );
  OAI222 U2396 ( .A(n1980), .B(n11038), .C(n1956), .D(n11271), .Q(n8832) );
  OAI222 U2397 ( .A(n1932), .B(n11036), .C(n1908), .D(n11270), .Q(n8831) );
  OAI222 U2399 ( .A(n2268), .B(n11034), .C(n2244), .D(n11269), .Q(n8838) );
  OAI222 U2400 ( .A(n2220), .B(n11032), .C(n2196), .D(n11268), .Q(n8837) );
  OAI222 U2401 ( .A(n2172), .B(n11030), .C(n2148), .D(n11267), .Q(n8836) );
  OAI222 U2402 ( .A(n2124), .B(n11028), .C(n2100), .D(n11266), .Q(n8835) );
  OAI222 U2405 ( .A(n924), .B(n11026), .C(n900), .D(n11265), .Q(n8846) );
  OAI222 U2406 ( .A(n876), .B(n11024), .C(n852), .D(n11264), .Q(n8845) );
  OAI222 U2407 ( .A(n828), .B(n11022), .C(n804), .D(n11263), .Q(n8844) );
  OAI222 U2408 ( .A(n780), .B(n11020), .C(n756), .D(n11262), .Q(n8843) );
  OAI222 U2410 ( .A(n1116), .B(n11018), .C(n1092), .D(n11261), .Q(n8850) );
  OAI222 U2411 ( .A(n1068), .B(n11016), .C(n1044), .D(n11260), .Q(n8849) );
  OAI222 U2412 ( .A(n1020), .B(n11014), .C(n996), .D(n11259), .Q(n8848) );
  OAI222 U2413 ( .A(n972), .B(n11012), .C(n948), .D(n11258), .Q(n8847) );
  OAI222 U2415 ( .A(n1308), .B(n11010), .C(n1284), .D(n11257), .Q(n8854) );
  OAI222 U2416 ( .A(n1260), .B(n11008), .C(n1236), .D(n11256), .Q(n8853) );
  OAI222 U2417 ( .A(n1212), .B(n11006), .C(n1188), .D(n11255), .Q(n8852) );
  OAI222 U2418 ( .A(n1164), .B(n11004), .C(n1140), .D(n11254), .Q(n8851) );
  OAI222 U2420 ( .A(n1500), .B(n11002), .C(n1476), .D(n11253), .Q(n8858) );
  OAI222 U2421 ( .A(n1452), .B(n11000), .C(n1428), .D(n11252), .Q(n8857) );
  OAI222 U2422 ( .A(n1404), .B(n10998), .C(n1380), .D(n11251), .Q(n8856) );
  OAI222 U2423 ( .A(n1356), .B(n10996), .C(n1332), .D(n11250), .Q(n8855) );
  OAI222 U2426 ( .A(n156), .B(n10994), .C(n132), .D(n11249), .Q(n8866) );
  OAI222 U2427 ( .A(n108), .B(n10992), .C(n84), .D(n11248), .Q(n8865) );
  OAI222 U2428 ( .A(n60), .B(n10990), .C(n36), .D(n11247), .Q(n8864) );
  OAI222 U2429 ( .A(n12), .B(n10988), .C(n6132), .D(n11246), .Q(n8863) );
  OAI222 U2431 ( .A(n348), .B(n10986), .C(n324), .D(n11245), .Q(n8870) );
  OAI222 U2432 ( .A(n300), .B(n10984), .C(n276), .D(n11244), .Q(n8869) );
  OAI222 U2433 ( .A(n252), .B(n10982), .C(n228), .D(n11243), .Q(n8868) );
  OAI222 U2434 ( .A(n204), .B(n10980), .C(n180), .D(n11242), .Q(n8867) );
  OAI222 U2436 ( .A(n540), .B(n10978), .C(n516), .D(n11241), .Q(n8874) );
  OAI222 U2437 ( .A(n492), .B(n10976), .C(n468), .D(n11240), .Q(n8873) );
  OAI222 U2438 ( .A(n444), .B(n10974), .C(n420), .D(n11239), .Q(n8872) );
  OAI222 U2439 ( .A(n396), .B(n10972), .C(n372), .D(n11238), .Q(n8871) );
  OAI222 U2441 ( .A(n732), .B(n10970), .C(n708), .D(n11237), .Q(n8878) );
  OAI222 U2442 ( .A(n684), .B(n10968), .C(n660), .D(n11236), .Q(n8877) );
  OAI222 U2443 ( .A(n636), .B(n10966), .C(n612), .D(n11235), .Q(n8876) );
  OAI222 U2444 ( .A(n588), .B(n10964), .C(n564), .D(n11234), .Q(n8875) );
  OAI222 U2448 ( .A(n5532), .B(n10962), .C(n5508), .D(n11233), .Q(n8890) );
  OAI222 U2449 ( .A(n5484), .B(n10960), .C(n5460), .D(n11232), .Q(n8889) );
  OAI222 U2450 ( .A(n5436), .B(n10958), .C(n5412), .D(n11231), .Q(n8888) );
  OAI222 U2451 ( .A(n5388), .B(n10956), .C(n5364), .D(n11230), .Q(n8887) );
  OAI222 U2453 ( .A(n5724), .B(n10954), .C(n5700), .D(n11229), .Q(n8894) );
  OAI222 U2454 ( .A(n5676), .B(n10952), .C(n5652), .D(n11228), .Q(n8893) );
  OAI222 U2455 ( .A(n5628), .B(n10950), .C(n5604), .D(n11227), .Q(n8892) );
  OAI222 U2456 ( .A(n5580), .B(n10948), .C(n5556), .D(n11226), .Q(n8891) );
  OAI222 U2458 ( .A(n5916), .B(n10946), .C(n5892), .D(n11225), .Q(n8898) );
  OAI222 U2459 ( .A(n5868), .B(n10944), .C(n5844), .D(n11224), .Q(n8897) );
  OAI222 U2460 ( .A(n5820), .B(n10942), .C(n5796), .D(n11223), .Q(n8896) );
  OAI222 U2461 ( .A(n5772), .B(n10940), .C(n5748), .D(n11222), .Q(n8895) );
  OAI222 U2463 ( .A(n6108), .B(n10938), .C(n6084), .D(n11221), .Q(n8902) );
  OAI222 U2464 ( .A(n6060), .B(n10936), .C(n6036), .D(n11220), .Q(n8901) );
  OAI222 U2465 ( .A(n6012), .B(n10934), .C(n5988), .D(n11219), .Q(n8900) );
  OAI222 U2466 ( .A(n5964), .B(n10932), .C(n5940), .D(n11218), .Q(n8899) );
  OAI222 U2469 ( .A(n4764), .B(n10930), .C(n4740), .D(n11217), .Q(n8910) );
  OAI222 U2470 ( .A(n4716), .B(n10928), .C(n4692), .D(n11216), .Q(n8909) );
  OAI222 U2471 ( .A(n4668), .B(n10926), .C(n4644), .D(n11215), .Q(n8908) );
  OAI222 U2472 ( .A(n4620), .B(n10924), .C(n4596), .D(n11214), .Q(n8907) );
  OAI222 U2474 ( .A(n4956), .B(n10922), .C(n4932), .D(n11213), .Q(n8914) );
  OAI222 U2475 ( .A(n4908), .B(n10920), .C(n4884), .D(n11212), .Q(n8913) );
  OAI222 U2476 ( .A(n4860), .B(n10918), .C(n4836), .D(n11211), .Q(n8912) );
  OAI222 U2477 ( .A(n4812), .B(n10916), .C(n4788), .D(n11210), .Q(n8911) );
  OAI222 U2479 ( .A(n5148), .B(n10914), .C(n5124), .D(n11209), .Q(n8918) );
  OAI222 U2480 ( .A(n5100), .B(n10912), .C(n5076), .D(n11208), .Q(n8917) );
  OAI222 U2481 ( .A(n5052), .B(n10910), .C(n5028), .D(n11207), .Q(n8916) );
  OAI222 U2482 ( .A(n5004), .B(n10908), .C(n4980), .D(n11206), .Q(n8915) );
  OAI222 U2484 ( .A(n5340), .B(n10906), .C(n5316), .D(n11205), .Q(n8922) );
  OAI222 U2485 ( .A(n5292), .B(n10904), .C(n5268), .D(n11204), .Q(n8921) );
  OAI222 U2486 ( .A(n5244), .B(n10902), .C(n5220), .D(n11203), .Q(n8920) );
  OAI222 U2487 ( .A(n5196), .B(n10900), .C(n5172), .D(n11202), .Q(n8919) );
  OAI222 U2490 ( .A(n3996), .B(n10898), .C(n3972), .D(n11201), .Q(n8930) );
  OAI222 U2491 ( .A(n3948), .B(n10896), .C(n3924), .D(n11200), .Q(n8929) );
  OAI222 U2492 ( .A(n3900), .B(n10894), .C(n3876), .D(n11199), .Q(n8928) );
  OAI222 U2493 ( .A(n3852), .B(n10892), .C(n3828), .D(n11198), .Q(n8927) );
  OAI222 U2495 ( .A(n4188), .B(n10890), .C(n4164), .D(n11197), .Q(n8934) );
  OAI222 U2496 ( .A(n4140), .B(n10888), .C(n4116), .D(n11196), .Q(n8933) );
  OAI222 U2497 ( .A(n4092), .B(n10886), .C(n4068), .D(n11195), .Q(n8932) );
  OAI222 U2498 ( .A(n4044), .B(n10884), .C(n4020), .D(n11194), .Q(n8931) );
  OAI222 U2500 ( .A(n4380), .B(n10882), .C(n4356), .D(n11193), .Q(n8938) );
  OAI222 U2501 ( .A(n4332), .B(n6192), .C(n4308), .D(n11192), .Q(n8937) );
  OAI222 U2502 ( .A(n4284), .B(n6190), .C(n4260), .D(n11191), .Q(n8936) );
  OAI222 U2503 ( .A(n4236), .B(n6188), .C(n4212), .D(n11190), .Q(n8935) );
  OAI222 U2505 ( .A(n4572), .B(n6186), .C(n4548), .D(n11189), .Q(n8942) );
  OAI222 U2506 ( .A(n4524), .B(n6184), .C(n4500), .D(n11188), .Q(n8941) );
  OAI222 U2507 ( .A(n4476), .B(n6182), .C(n4452), .D(n11187), .Q(n8940) );
  OAI222 U2508 ( .A(n4428), .B(n6180), .C(n4404), .D(n11186), .Q(n8939) );
  OAI222 U2511 ( .A(n3228), .B(n6178), .C(n3204), .D(n11185), .Q(n8950) );
  OAI222 U2512 ( .A(n3180), .B(n6176), .C(n3156), .D(n11184), .Q(n8949) );
  OAI222 U2513 ( .A(n3132), .B(n6174), .C(n3108), .D(n11183), .Q(n8948) );
  OAI222 U2514 ( .A(n3084), .B(n6172), .C(n3060), .D(n11182), .Q(n8947) );
  OAI222 U2516 ( .A(n3420), .B(n6170), .C(n3396), .D(n11181), .Q(n8954) );
  OAI222 U2517 ( .A(n3372), .B(n6168), .C(n3348), .D(n11180), .Q(n8953) );
  OAI222 U2518 ( .A(n3324), .B(n6166), .C(n3300), .D(n11179), .Q(n8952) );
  OAI222 U2519 ( .A(n3276), .B(n6164), .C(n3252), .D(n11178), .Q(n8951) );
  OAI222 U2521 ( .A(n3612), .B(n6162), .C(n3588), .D(n11177), .Q(n8958) );
  OAI222 U2522 ( .A(n3564), .B(n6160), .C(n3540), .D(n11176), .Q(n8957) );
  OAI222 U2523 ( .A(n3516), .B(n6158), .C(n3492), .D(n11175), .Q(n8956) );
  OAI222 U2524 ( .A(n3468), .B(n6156), .C(n3444), .D(n11174), .Q(n8955) );
  OAI222 U2526 ( .A(n3804), .B(n6154), .C(n3780), .D(n11173), .Q(n8962) );
  OAI222 U2527 ( .A(n3756), .B(n6152), .C(n3732), .D(n11172), .Q(n8961) );
  OAI222 U2528 ( .A(n3708), .B(n6150), .C(n3684), .D(n11171), .Q(n8960) );
  OAI222 U2529 ( .A(n3660), .B(n6148), .C(n3636), .D(n11170), .Q(n8959) );
  OAI222 U2534 ( .A(n2459), .B(n11090), .C(n2435), .D(n11297), .Q(n8976) );
  OAI222 U2535 ( .A(n2411), .B(n11088), .C(n2387), .D(n11296), .Q(n8975) );
  OAI222 U2536 ( .A(n2363), .B(n11086), .C(n2339), .D(n11295), .Q(n8974) );
  OAI222 U2537 ( .A(n2315), .B(n11084), .C(n2291), .D(n11294), .Q(n8973) );
  OAI222 U2539 ( .A(n2651), .B(n11082), .C(n2627), .D(n11293), .Q(n8980) );
  OAI222 U2540 ( .A(n2603), .B(n11080), .C(n2579), .D(n11292), .Q(n8979) );
  OAI222 U2541 ( .A(n2555), .B(n11078), .C(n2531), .D(n11291), .Q(n8978) );
  OAI222 U2542 ( .A(n2507), .B(n11076), .C(n2483), .D(n11290), .Q(n8977) );
  OAI222 U2544 ( .A(n2843), .B(n11074), .C(n2819), .D(n11289), .Q(n8984) );
  OAI222 U2545 ( .A(n2795), .B(n11072), .C(n2771), .D(n11288), .Q(n8983) );
  OAI222 U2546 ( .A(n2747), .B(n11070), .C(n2723), .D(n11287), .Q(n8982) );
  OAI222 U2547 ( .A(n2699), .B(n11068), .C(n2675), .D(n11286), .Q(n8981) );
  OAI222 U2549 ( .A(n3035), .B(n11066), .C(n3011), .D(n11285), .Q(n8988) );
  OAI222 U2550 ( .A(n2987), .B(n11064), .C(n2963), .D(n11284), .Q(n8987) );
  OAI222 U2551 ( .A(n2939), .B(n11062), .C(n2915), .D(n11283), .Q(n8986) );
  OAI222 U2552 ( .A(n2891), .B(n11060), .C(n2867), .D(n11282), .Q(n8985) );
  OAI222 U2555 ( .A(n1691), .B(n11058), .C(n1667), .D(n11281), .Q(n8996) );
  OAI222 U2556 ( .A(n1643), .B(n11056), .C(n1619), .D(n11280), .Q(n8995) );
  OAI222 U2557 ( .A(n1595), .B(n11054), .C(n1571), .D(n11279), .Q(n8994) );
  OAI222 U2558 ( .A(n1547), .B(n11052), .C(n1523), .D(n11278), .Q(n8993) );
  OAI222 U2560 ( .A(n1883), .B(n11050), .C(n1859), .D(n11277), .Q(n9000) );
  OAI222 U2561 ( .A(n1835), .B(n11048), .C(n1811), .D(n11276), .Q(n8999) );
  OAI222 U2562 ( .A(n1787), .B(n11046), .C(n1763), .D(n11275), .Q(n8998) );
  OAI222 U2563 ( .A(n1739), .B(n11044), .C(n1715), .D(n11274), .Q(n8997) );
  OAI222 U2565 ( .A(n2075), .B(n11042), .C(n2051), .D(n11273), .Q(n9004) );
  OAI222 U2566 ( .A(n2027), .B(n11040), .C(n2003), .D(n11272), .Q(n9003) );
  OAI222 U2567 ( .A(n1979), .B(n11038), .C(n1955), .D(n11271), .Q(n9002) );
  OAI222 U2568 ( .A(n1931), .B(n11036), .C(n1907), .D(n11270), .Q(n9001) );
  OAI222 U2570 ( .A(n2267), .B(n11034), .C(n2243), .D(n11269), .Q(n9008) );
  OAI222 U2571 ( .A(n2219), .B(n11032), .C(n2195), .D(n11268), .Q(n9007) );
  OAI222 U2572 ( .A(n2171), .B(n11030), .C(n2147), .D(n11267), .Q(n9006) );
  OAI222 U2573 ( .A(n2123), .B(n11028), .C(n2099), .D(n11266), .Q(n9005) );
  OAI222 U2576 ( .A(n923), .B(n11026), .C(n899), .D(n11265), .Q(n9016) );
  OAI222 U2577 ( .A(n875), .B(n11024), .C(n851), .D(n11264), .Q(n9015) );
  OAI222 U2578 ( .A(n827), .B(n11022), .C(n803), .D(n11263), .Q(n9014) );
  OAI222 U2579 ( .A(n779), .B(n11020), .C(n755), .D(n11262), .Q(n9013) );
  OAI222 U2581 ( .A(n1115), .B(n11018), .C(n1091), .D(n11261), .Q(n9020) );
  OAI222 U2582 ( .A(n1067), .B(n11016), .C(n1043), .D(n11260), .Q(n9019) );
  OAI222 U2583 ( .A(n1019), .B(n11014), .C(n995), .D(n11259), .Q(n9018) );
  OAI222 U2584 ( .A(n971), .B(n11012), .C(n947), .D(n11258), .Q(n9017) );
  OAI222 U2586 ( .A(n1307), .B(n11010), .C(n1283), .D(n11257), .Q(n9024) );
  OAI222 U2587 ( .A(n1259), .B(n11008), .C(n1235), .D(n11256), .Q(n9023) );
  OAI222 U2588 ( .A(n1211), .B(n11006), .C(n1187), .D(n11255), .Q(n9022) );
  OAI222 U2589 ( .A(n1163), .B(n11004), .C(n1139), .D(n11254), .Q(n9021) );
  OAI222 U2591 ( .A(n1499), .B(n11002), .C(n1475), .D(n11253), .Q(n9028) );
  OAI222 U2592 ( .A(n1451), .B(n11000), .C(n1427), .D(n11252), .Q(n9027) );
  OAI222 U2593 ( .A(n1403), .B(n10998), .C(n1379), .D(n11251), .Q(n9026) );
  OAI222 U2594 ( .A(n1355), .B(n10996), .C(n1331), .D(n11250), .Q(n9025) );
  OAI222 U2597 ( .A(n155), .B(n10994), .C(n131), .D(n11249), .Q(n9036) );
  OAI222 U2598 ( .A(n107), .B(n10992), .C(n83), .D(n11248), .Q(n9035) );
  OAI222 U2599 ( .A(n59), .B(n10990), .C(n35), .D(n11247), .Q(n9034) );
  OAI222 U2600 ( .A(n11), .B(n10988), .C(n6131), .D(n11246), .Q(n9033) );
  OAI222 U2602 ( .A(n347), .B(n10986), .C(n323), .D(n11245), .Q(n9040) );
  OAI222 U2603 ( .A(n299), .B(n10984), .C(n275), .D(n11244), .Q(n9039) );
  OAI222 U2604 ( .A(n251), .B(n10982), .C(n227), .D(n11243), .Q(n9038) );
  OAI222 U2605 ( .A(n203), .B(n10980), .C(n179), .D(n11242), .Q(n9037) );
  OAI222 U2607 ( .A(n539), .B(n10978), .C(n515), .D(n11241), .Q(n9044) );
  OAI222 U2608 ( .A(n491), .B(n10976), .C(n467), .D(n11240), .Q(n9043) );
  OAI222 U2609 ( .A(n443), .B(n10974), .C(n419), .D(n11239), .Q(n9042) );
  OAI222 U2610 ( .A(n395), .B(n10972), .C(n371), .D(n11238), .Q(n9041) );
  OAI222 U2612 ( .A(n731), .B(n10970), .C(n707), .D(n11237), .Q(n9048) );
  OAI222 U2613 ( .A(n683), .B(n10968), .C(n659), .D(n11236), .Q(n9047) );
  OAI222 U2614 ( .A(n635), .B(n10966), .C(n611), .D(n11235), .Q(n9046) );
  OAI222 U2615 ( .A(n587), .B(n10964), .C(n563), .D(n11234), .Q(n9045) );
  OAI222 U2619 ( .A(n5531), .B(n10962), .C(n5507), .D(n11233), .Q(n9060) );
  OAI222 U2620 ( .A(n5483), .B(n10960), .C(n5459), .D(n11232), .Q(n9059) );
  OAI222 U2621 ( .A(n5435), .B(n10958), .C(n5411), .D(n11231), .Q(n9058) );
  OAI222 U2622 ( .A(n5387), .B(n10956), .C(n5363), .D(n11230), .Q(n9057) );
  OAI222 U2624 ( .A(n5723), .B(n10954), .C(n5699), .D(n11229), .Q(n9064) );
  OAI222 U2625 ( .A(n5675), .B(n10952), .C(n5651), .D(n11228), .Q(n9063) );
  OAI222 U2626 ( .A(n5627), .B(n10950), .C(n5603), .D(n11227), .Q(n9062) );
  OAI222 U2627 ( .A(n5579), .B(n10948), .C(n5555), .D(n11226), .Q(n9061) );
  OAI222 U2629 ( .A(n5915), .B(n10946), .C(n5891), .D(n11225), .Q(n9068) );
  OAI222 U2630 ( .A(n5867), .B(n10944), .C(n5843), .D(n11224), .Q(n9067) );
  OAI222 U2631 ( .A(n5819), .B(n10942), .C(n5795), .D(n11223), .Q(n9066) );
  OAI222 U2632 ( .A(n5771), .B(n10940), .C(n5747), .D(n11222), .Q(n9065) );
  OAI222 U2634 ( .A(n6107), .B(n10938), .C(n6083), .D(n11221), .Q(n9072) );
  OAI222 U2635 ( .A(n6059), .B(n10936), .C(n6035), .D(n11220), .Q(n9071) );
  OAI222 U2636 ( .A(n6011), .B(n10934), .C(n5987), .D(n11219), .Q(n9070) );
  OAI222 U2637 ( .A(n5963), .B(n10932), .C(n5939), .D(n11218), .Q(n9069) );
  OAI222 U2640 ( .A(n4763), .B(n10930), .C(n4739), .D(n11217), .Q(n9080) );
  OAI222 U2641 ( .A(n4715), .B(n10928), .C(n4691), .D(n11216), .Q(n9079) );
  OAI222 U2642 ( .A(n4667), .B(n10926), .C(n4643), .D(n11215), .Q(n9078) );
  OAI222 U2643 ( .A(n4619), .B(n10924), .C(n4595), .D(n11214), .Q(n9077) );
  OAI222 U2645 ( .A(n4955), .B(n10922), .C(n4931), .D(n11213), .Q(n9084) );
  OAI222 U2646 ( .A(n4907), .B(n10920), .C(n4883), .D(n11212), .Q(n9083) );
  OAI222 U2647 ( .A(n4859), .B(n10918), .C(n4835), .D(n11211), .Q(n9082) );
  OAI222 U2648 ( .A(n4811), .B(n10916), .C(n4787), .D(n11210), .Q(n9081) );
  OAI222 U2650 ( .A(n5147), .B(n10914), .C(n5123), .D(n11209), .Q(n9088) );
  OAI222 U2651 ( .A(n5099), .B(n10912), .C(n5075), .D(n11208), .Q(n9087) );
  OAI222 U2652 ( .A(n5051), .B(n10910), .C(n5027), .D(n11207), .Q(n9086) );
  OAI222 U2653 ( .A(n5003), .B(n10908), .C(n4979), .D(n11206), .Q(n9085) );
  OAI222 U2655 ( .A(n5339), .B(n10906), .C(n5315), .D(n11205), .Q(n9092) );
  OAI222 U2656 ( .A(n5291), .B(n10904), .C(n5267), .D(n11204), .Q(n9091) );
  OAI222 U2657 ( .A(n5243), .B(n10902), .C(n5219), .D(n11203), .Q(n9090) );
  OAI222 U2658 ( .A(n5195), .B(n10900), .C(n5171), .D(n11202), .Q(n9089) );
  OAI222 U2661 ( .A(n3995), .B(n10898), .C(n3971), .D(n11201), .Q(n9100) );
  OAI222 U2662 ( .A(n3947), .B(n10896), .C(n3923), .D(n11200), .Q(n9099) );
  OAI222 U2663 ( .A(n3899), .B(n10894), .C(n3875), .D(n11199), .Q(n9098) );
  OAI222 U2664 ( .A(n3851), .B(n10892), .C(n3827), .D(n11198), .Q(n9097) );
  OAI222 U2666 ( .A(n4187), .B(n10890), .C(n4163), .D(n11197), .Q(n9104) );
  OAI222 U2667 ( .A(n4139), .B(n10888), .C(n4115), .D(n11196), .Q(n9103) );
  OAI222 U2668 ( .A(n4091), .B(n10886), .C(n4067), .D(n11195), .Q(n9102) );
  OAI222 U2669 ( .A(n4043), .B(n10884), .C(n4019), .D(n11194), .Q(n9101) );
  OAI222 U2671 ( .A(n4379), .B(n10882), .C(n4355), .D(n11193), .Q(n9108) );
  OAI222 U2672 ( .A(n4331), .B(n6192), .C(n4307), .D(n11192), .Q(n9107) );
  OAI222 U2673 ( .A(n4283), .B(n6190), .C(n4259), .D(n11191), .Q(n9106) );
  OAI222 U2674 ( .A(n4235), .B(n6188), .C(n4211), .D(n11190), .Q(n9105) );
  OAI222 U2676 ( .A(n4571), .B(n6186), .C(n4547), .D(n11189), .Q(n9112) );
  OAI222 U2677 ( .A(n4523), .B(n6184), .C(n4499), .D(n11188), .Q(n9111) );
  OAI222 U2678 ( .A(n4475), .B(n6182), .C(n4451), .D(n11187), .Q(n9110) );
  OAI222 U2679 ( .A(n4427), .B(n6180), .C(n4403), .D(n11186), .Q(n9109) );
  OAI222 U2682 ( .A(n3227), .B(n6178), .C(n3203), .D(n11185), .Q(n9120) );
  OAI222 U2683 ( .A(n3179), .B(n6176), .C(n3155), .D(n11184), .Q(n9119) );
  OAI222 U2684 ( .A(n3131), .B(n6174), .C(n3107), .D(n11183), .Q(n9118) );
  OAI222 U2685 ( .A(n3083), .B(n6172), .C(n3059), .D(n11182), .Q(n9117) );
  OAI222 U2687 ( .A(n3419), .B(n6170), .C(n3395), .D(n11181), .Q(n9124) );
  OAI222 U2688 ( .A(n3371), .B(n6168), .C(n3347), .D(n11180), .Q(n9123) );
  OAI222 U2689 ( .A(n3323), .B(n6166), .C(n3299), .D(n11179), .Q(n9122) );
  OAI222 U2690 ( .A(n3275), .B(n6164), .C(n3251), .D(n11178), .Q(n9121) );
  OAI222 U2692 ( .A(n3611), .B(n6162), .C(n3587), .D(n11177), .Q(n9128) );
  OAI222 U2693 ( .A(n3563), .B(n6160), .C(n3539), .D(n11176), .Q(n9127) );
  OAI222 U2694 ( .A(n3515), .B(n6158), .C(n3491), .D(n11175), .Q(n9126) );
  OAI222 U2695 ( .A(n3467), .B(n6156), .C(n3443), .D(n11174), .Q(n9125) );
  OAI222 U2697 ( .A(n3803), .B(n6154), .C(n3779), .D(n11173), .Q(n9132) );
  OAI222 U2698 ( .A(n3755), .B(n6152), .C(n3731), .D(n11172), .Q(n9131) );
  OAI222 U2699 ( .A(n3707), .B(n6150), .C(n3683), .D(n11171), .Q(n9130) );
  OAI222 U2700 ( .A(n3659), .B(n6148), .C(n3635), .D(n11170), .Q(n9129) );
  OAI222 U2705 ( .A(n2458), .B(n11090), .C(n2434), .D(n11297), .Q(n9146) );
  OAI222 U2706 ( .A(n2410), .B(n11088), .C(n2386), .D(n11296), .Q(n9145) );
  OAI222 U2707 ( .A(n2362), .B(n11086), .C(n2338), .D(n11295), .Q(n9144) );
  OAI222 U2708 ( .A(n2314), .B(n11084), .C(n2290), .D(n11294), .Q(n9143) );
  OAI222 U2710 ( .A(n2650), .B(n11082), .C(n2626), .D(n11293), .Q(n9150) );
  OAI222 U2711 ( .A(n2602), .B(n11080), .C(n2578), .D(n11292), .Q(n9149) );
  OAI222 U2712 ( .A(n2554), .B(n11078), .C(n2530), .D(n11291), .Q(n9148) );
  OAI222 U2713 ( .A(n2506), .B(n11076), .C(n2482), .D(n11290), .Q(n9147) );
  OAI222 U2715 ( .A(n2842), .B(n11074), .C(n2818), .D(n11289), .Q(n9154) );
  OAI222 U2716 ( .A(n2794), .B(n11072), .C(n2770), .D(n11288), .Q(n9153) );
  OAI222 U2717 ( .A(n2746), .B(n11070), .C(n2722), .D(n11287), .Q(n9152) );
  OAI222 U2718 ( .A(n2698), .B(n11068), .C(n2674), .D(n11286), .Q(n9151) );
  OAI222 U2720 ( .A(n3034), .B(n11066), .C(n3010), .D(n11285), .Q(n9158) );
  OAI222 U2721 ( .A(n2986), .B(n11064), .C(n2962), .D(n11284), .Q(n9157) );
  OAI222 U2722 ( .A(n2938), .B(n11062), .C(n2914), .D(n11283), .Q(n9156) );
  OAI222 U2723 ( .A(n2890), .B(n11060), .C(n2866), .D(n11282), .Q(n9155) );
  OAI222 U2726 ( .A(n1690), .B(n11058), .C(n1666), .D(n11281), .Q(n9166) );
  OAI222 U2727 ( .A(n1642), .B(n11056), .C(n1618), .D(n11280), .Q(n9165) );
  OAI222 U2728 ( .A(n1594), .B(n11054), .C(n1570), .D(n11279), .Q(n9164) );
  OAI222 U2729 ( .A(n1546), .B(n11052), .C(n1522), .D(n11278), .Q(n9163) );
  OAI222 U2731 ( .A(n1882), .B(n11050), .C(n1858), .D(n11277), .Q(n9170) );
  OAI222 U2732 ( .A(n1834), .B(n11048), .C(n1810), .D(n11276), .Q(n9169) );
  OAI222 U2733 ( .A(n1786), .B(n11046), .C(n1762), .D(n11275), .Q(n9168) );
  OAI222 U2734 ( .A(n1738), .B(n11044), .C(n1714), .D(n11274), .Q(n9167) );
  OAI222 U2736 ( .A(n2074), .B(n11042), .C(n2050), .D(n11273), .Q(n9174) );
  OAI222 U2737 ( .A(n2026), .B(n11040), .C(n2002), .D(n11272), .Q(n9173) );
  OAI222 U2738 ( .A(n1978), .B(n11038), .C(n1954), .D(n11271), .Q(n9172) );
  OAI222 U2739 ( .A(n1930), .B(n11036), .C(n1906), .D(n11270), .Q(n9171) );
  OAI222 U2741 ( .A(n2266), .B(n11034), .C(n2242), .D(n11269), .Q(n9178) );
  OAI222 U2742 ( .A(n2218), .B(n11032), .C(n2194), .D(n11268), .Q(n9177) );
  OAI222 U2743 ( .A(n2170), .B(n11030), .C(n2146), .D(n11267), .Q(n9176) );
  OAI222 U2744 ( .A(n2122), .B(n11028), .C(n2098), .D(n11266), .Q(n9175) );
  OAI222 U2747 ( .A(n922), .B(n11026), .C(n898), .D(n11265), .Q(n9186) );
  OAI222 U2748 ( .A(n874), .B(n11024), .C(n850), .D(n11264), .Q(n9185) );
  OAI222 U2749 ( .A(n826), .B(n11022), .C(n802), .D(n11263), .Q(n9184) );
  OAI222 U2750 ( .A(n778), .B(n11020), .C(n754), .D(n11262), .Q(n9183) );
  OAI222 U2752 ( .A(n1114), .B(n11018), .C(n1090), .D(n11261), .Q(n9190) );
  OAI222 U2753 ( .A(n1066), .B(n11016), .C(n1042), .D(n11260), .Q(n9189) );
  OAI222 U2754 ( .A(n1018), .B(n11014), .C(n994), .D(n11259), .Q(n9188) );
  OAI222 U2755 ( .A(n970), .B(n11012), .C(n946), .D(n11258), .Q(n9187) );
  OAI222 U2757 ( .A(n1306), .B(n11010), .C(n1282), .D(n11257), .Q(n9194) );
  OAI222 U2758 ( .A(n1258), .B(n11008), .C(n1234), .D(n11256), .Q(n9193) );
  OAI222 U2759 ( .A(n1210), .B(n11006), .C(n1186), .D(n11255), .Q(n9192) );
  OAI222 U2760 ( .A(n1162), .B(n11004), .C(n1138), .D(n11254), .Q(n9191) );
  OAI222 U2762 ( .A(n1498), .B(n11002), .C(n1474), .D(n11253), .Q(n9198) );
  OAI222 U2763 ( .A(n1450), .B(n11000), .C(n1426), .D(n11252), .Q(n9197) );
  OAI222 U2764 ( .A(n1402), .B(n10998), .C(n1378), .D(n11251), .Q(n9196) );
  OAI222 U2765 ( .A(n1354), .B(n10996), .C(n1330), .D(n11250), .Q(n9195) );
  OAI222 U2768 ( .A(n154), .B(n10994), .C(n130), .D(n11249), .Q(n9206) );
  OAI222 U2769 ( .A(n106), .B(n10992), .C(n82), .D(n11248), .Q(n9205) );
  OAI222 U2770 ( .A(n58), .B(n10990), .C(n34), .D(n11247), .Q(n9204) );
  OAI222 U2771 ( .A(n10), .B(n10988), .C(n6130), .D(n11246), .Q(n9203) );
  OAI222 U2773 ( .A(n346), .B(n10986), .C(n322), .D(n11245), .Q(n9210) );
  OAI222 U2774 ( .A(n298), .B(n10984), .C(n274), .D(n11244), .Q(n9209) );
  OAI222 U2775 ( .A(n250), .B(n10982), .C(n226), .D(n11243), .Q(n9208) );
  OAI222 U2776 ( .A(n202), .B(n10980), .C(n178), .D(n11242), .Q(n9207) );
  OAI222 U2778 ( .A(n538), .B(n10978), .C(n514), .D(n11241), .Q(n9214) );
  OAI222 U2779 ( .A(n490), .B(n10976), .C(n466), .D(n11240), .Q(n9213) );
  OAI222 U2780 ( .A(n442), .B(n10974), .C(n418), .D(n11239), .Q(n9212) );
  OAI222 U2781 ( .A(n394), .B(n10972), .C(n370), .D(n11238), .Q(n9211) );
  OAI222 U2783 ( .A(n730), .B(n10970), .C(n706), .D(n11237), .Q(n9218) );
  OAI222 U2784 ( .A(n682), .B(n10968), .C(n658), .D(n11236), .Q(n9217) );
  OAI222 U2785 ( .A(n634), .B(n10966), .C(n610), .D(n11235), .Q(n9216) );
  OAI222 U2786 ( .A(n586), .B(n10964), .C(n562), .D(n11234), .Q(n9215) );
  OAI222 U2790 ( .A(n5530), .B(n10962), .C(n5506), .D(n11233), .Q(n9230) );
  OAI222 U2791 ( .A(n5482), .B(n10960), .C(n5458), .D(n11232), .Q(n9229) );
  OAI222 U2792 ( .A(n5434), .B(n10958), .C(n5410), .D(n11231), .Q(n9228) );
  OAI222 U2793 ( .A(n5386), .B(n10956), .C(n5362), .D(n11230), .Q(n9227) );
  OAI222 U2795 ( .A(n5722), .B(n10954), .C(n5698), .D(n11229), .Q(n9234) );
  OAI222 U2796 ( .A(n5674), .B(n10952), .C(n5650), .D(n11228), .Q(n9233) );
  OAI222 U2797 ( .A(n5626), .B(n10950), .C(n5602), .D(n11227), .Q(n9232) );
  OAI222 U2798 ( .A(n5578), .B(n10948), .C(n5554), .D(n11226), .Q(n9231) );
  OAI222 U2800 ( .A(n5914), .B(n10946), .C(n5890), .D(n11225), .Q(n9238) );
  OAI222 U2801 ( .A(n5866), .B(n10944), .C(n5842), .D(n11224), .Q(n9237) );
  OAI222 U2802 ( .A(n5818), .B(n10942), .C(n5794), .D(n11223), .Q(n9236) );
  OAI222 U2803 ( .A(n5770), .B(n10940), .C(n5746), .D(n11222), .Q(n9235) );
  OAI222 U2805 ( .A(n6106), .B(n10938), .C(n6082), .D(n11221), .Q(n9242) );
  OAI222 U2806 ( .A(n6058), .B(n10936), .C(n6034), .D(n11220), .Q(n9241) );
  OAI222 U2807 ( .A(n6010), .B(n10934), .C(n5986), .D(n11219), .Q(n9240) );
  OAI222 U2808 ( .A(n5962), .B(n10932), .C(n5938), .D(n11218), .Q(n9239) );
  OAI222 U2811 ( .A(n4762), .B(n10930), .C(n4738), .D(n11217), .Q(n9250) );
  OAI222 U2812 ( .A(n4714), .B(n10928), .C(n4690), .D(n11216), .Q(n9249) );
  OAI222 U2813 ( .A(n4666), .B(n10926), .C(n4642), .D(n11215), .Q(n9248) );
  OAI222 U2814 ( .A(n4618), .B(n10924), .C(n4594), .D(n11214), .Q(n9247) );
  OAI222 U2816 ( .A(n4954), .B(n10922), .C(n4930), .D(n11213), .Q(n9254) );
  OAI222 U2817 ( .A(n4906), .B(n10920), .C(n4882), .D(n11212), .Q(n9253) );
  OAI222 U2818 ( .A(n4858), .B(n10918), .C(n4834), .D(n11211), .Q(n9252) );
  OAI222 U2819 ( .A(n4810), .B(n10916), .C(n4786), .D(n11210), .Q(n9251) );
  OAI222 U2821 ( .A(n5146), .B(n10914), .C(n5122), .D(n11209), .Q(n9258) );
  OAI222 U2822 ( .A(n5098), .B(n10912), .C(n5074), .D(n11208), .Q(n9257) );
  OAI222 U2823 ( .A(n5050), .B(n10910), .C(n5026), .D(n11207), .Q(n9256) );
  OAI222 U2824 ( .A(n5002), .B(n10908), .C(n4978), .D(n11206), .Q(n9255) );
  OAI222 U2826 ( .A(n5338), .B(n10906), .C(n5314), .D(n11205), .Q(n9262) );
  OAI222 U2827 ( .A(n5290), .B(n10904), .C(n5266), .D(n11204), .Q(n9261) );
  OAI222 U2828 ( .A(n5242), .B(n10902), .C(n5218), .D(n11203), .Q(n9260) );
  OAI222 U2829 ( .A(n5194), .B(n10900), .C(n5170), .D(n11202), .Q(n9259) );
  OAI222 U2832 ( .A(n3994), .B(n10898), .C(n3970), .D(n11201), .Q(n9270) );
  OAI222 U2833 ( .A(n3946), .B(n10896), .C(n3922), .D(n11200), .Q(n9269) );
  OAI222 U2834 ( .A(n3898), .B(n10894), .C(n3874), .D(n11199), .Q(n9268) );
  OAI222 U2835 ( .A(n3850), .B(n10892), .C(n3826), .D(n11198), .Q(n9267) );
  OAI222 U2837 ( .A(n4186), .B(n10890), .C(n4162), .D(n11197), .Q(n9274) );
  OAI222 U2838 ( .A(n4138), .B(n10888), .C(n4114), .D(n11196), .Q(n9273) );
  OAI222 U2839 ( .A(n4090), .B(n10886), .C(n4066), .D(n11195), .Q(n9272) );
  OAI222 U2840 ( .A(n4042), .B(n10884), .C(n4018), .D(n11194), .Q(n9271) );
  OAI222 U2842 ( .A(n4378), .B(n10882), .C(n4354), .D(n11193), .Q(n9278) );
  OAI222 U2843 ( .A(n4330), .B(n6192), .C(n4306), .D(n11192), .Q(n9277) );
  OAI222 U2844 ( .A(n4282), .B(n6190), .C(n4258), .D(n11191), .Q(n9276) );
  OAI222 U2845 ( .A(n4234), .B(n6188), .C(n4210), .D(n11190), .Q(n9275) );
  OAI222 U2847 ( .A(n4570), .B(n6186), .C(n4546), .D(n11189), .Q(n9282) );
  OAI222 U2848 ( .A(n4522), .B(n6184), .C(n4498), .D(n11188), .Q(n9281) );
  OAI222 U2849 ( .A(n4474), .B(n6182), .C(n4450), .D(n11187), .Q(n9280) );
  OAI222 U2850 ( .A(n4426), .B(n6180), .C(n4402), .D(n11186), .Q(n9279) );
  OAI222 U2853 ( .A(n3226), .B(n6178), .C(n3202), .D(n11185), .Q(n9290) );
  OAI222 U2854 ( .A(n3178), .B(n6176), .C(n3154), .D(n11184), .Q(n9289) );
  OAI222 U2855 ( .A(n3130), .B(n6174), .C(n3106), .D(n11183), .Q(n9288) );
  OAI222 U2856 ( .A(n3082), .B(n6172), .C(n3058), .D(n11182), .Q(n9287) );
  OAI222 U2858 ( .A(n3418), .B(n6170), .C(n3394), .D(n11181), .Q(n9294) );
  OAI222 U2859 ( .A(n3370), .B(n6168), .C(n3346), .D(n11180), .Q(n9293) );
  OAI222 U2860 ( .A(n3322), .B(n6166), .C(n3298), .D(n11179), .Q(n9292) );
  OAI222 U2861 ( .A(n3274), .B(n6164), .C(n3250), .D(n11178), .Q(n9291) );
  OAI222 U2863 ( .A(n3610), .B(n6162), .C(n3586), .D(n11177), .Q(n9298) );
  OAI222 U2864 ( .A(n3562), .B(n6160), .C(n3538), .D(n11176), .Q(n9297) );
  OAI222 U2865 ( .A(n3514), .B(n6158), .C(n3490), .D(n11175), .Q(n9296) );
  OAI222 U2866 ( .A(n3466), .B(n6156), .C(n3442), .D(n11174), .Q(n9295) );
  OAI222 U2868 ( .A(n3802), .B(n6154), .C(n3778), .D(n11173), .Q(n9302) );
  OAI222 U2869 ( .A(n3754), .B(n6152), .C(n3730), .D(n11172), .Q(n9301) );
  OAI222 U2870 ( .A(n3706), .B(n6150), .C(n3682), .D(n11171), .Q(n9300) );
  OAI222 U2871 ( .A(n3658), .B(n6148), .C(n3634), .D(n11170), .Q(n9299) );
  OAI222 U2876 ( .A(n2457), .B(n11090), .C(n2433), .D(n11297), .Q(n9316) );
  OAI222 U2877 ( .A(n2409), .B(n11088), .C(n2385), .D(n11296), .Q(n9315) );
  OAI222 U2878 ( .A(n2361), .B(n11086), .C(n2337), .D(n11295), .Q(n9314) );
  OAI222 U2879 ( .A(n2313), .B(n11084), .C(n2289), .D(n11294), .Q(n9313) );
  OAI222 U2881 ( .A(n2649), .B(n11082), .C(n2625), .D(n11293), .Q(n9320) );
  OAI222 U2882 ( .A(n2601), .B(n11080), .C(n2577), .D(n11292), .Q(n9319) );
  OAI222 U2883 ( .A(n2553), .B(n11078), .C(n2529), .D(n11291), .Q(n9318) );
  OAI222 U2884 ( .A(n2505), .B(n11076), .C(n2481), .D(n11290), .Q(n9317) );
  OAI222 U2886 ( .A(n2841), .B(n11074), .C(n2817), .D(n11289), .Q(n9324) );
  OAI222 U2887 ( .A(n2793), .B(n11072), .C(n2769), .D(n11288), .Q(n9323) );
  OAI222 U2888 ( .A(n2745), .B(n11070), .C(n2721), .D(n11287), .Q(n9322) );
  OAI222 U2889 ( .A(n2697), .B(n11068), .C(n2673), .D(n11286), .Q(n9321) );
  OAI222 U2891 ( .A(n3033), .B(n11066), .C(n3009), .D(n11285), .Q(n9328) );
  OAI222 U2892 ( .A(n2985), .B(n11064), .C(n2961), .D(n11284), .Q(n9327) );
  OAI222 U2893 ( .A(n2937), .B(n11062), .C(n2913), .D(n11283), .Q(n9326) );
  OAI222 U2894 ( .A(n2889), .B(n11060), .C(n2865), .D(n11282), .Q(n9325) );
  OAI222 U2897 ( .A(n1689), .B(n11058), .C(n1665), .D(n11281), .Q(n9336) );
  OAI222 U2898 ( .A(n1641), .B(n11056), .C(n1617), .D(n11280), .Q(n9335) );
  OAI222 U2899 ( .A(n1593), .B(n11054), .C(n1569), .D(n11279), .Q(n9334) );
  OAI222 U2900 ( .A(n1545), .B(n11052), .C(n1521), .D(n11278), .Q(n9333) );
  OAI222 U2902 ( .A(n1881), .B(n11050), .C(n1857), .D(n11277), .Q(n9340) );
  OAI222 U2903 ( .A(n1833), .B(n11048), .C(n1809), .D(n11276), .Q(n9339) );
  OAI222 U2904 ( .A(n1785), .B(n11046), .C(n1761), .D(n11275), .Q(n9338) );
  OAI222 U2905 ( .A(n1737), .B(n11044), .C(n1713), .D(n11274), .Q(n9337) );
  OAI222 U2907 ( .A(n2073), .B(n11042), .C(n2049), .D(n11273), .Q(n9344) );
  OAI222 U2908 ( .A(n2025), .B(n11040), .C(n2001), .D(n11272), .Q(n9343) );
  OAI222 U2909 ( .A(n1977), .B(n11038), .C(n1953), .D(n11271), .Q(n9342) );
  OAI222 U2910 ( .A(n1929), .B(n11036), .C(n1905), .D(n11270), .Q(n9341) );
  OAI222 U2912 ( .A(n2265), .B(n11034), .C(n2241), .D(n11269), .Q(n9348) );
  OAI222 U2913 ( .A(n2217), .B(n11032), .C(n2193), .D(n11268), .Q(n9347) );
  OAI222 U2914 ( .A(n2169), .B(n11030), .C(n2145), .D(n11267), .Q(n9346) );
  OAI222 U2915 ( .A(n2121), .B(n11028), .C(n2097), .D(n11266), .Q(n9345) );
  OAI222 U2918 ( .A(n921), .B(n11026), .C(n897), .D(n11265), .Q(n9356) );
  OAI222 U2919 ( .A(n873), .B(n11024), .C(n849), .D(n11264), .Q(n9355) );
  OAI222 U2920 ( .A(n825), .B(n11022), .C(n801), .D(n11263), .Q(n9354) );
  OAI222 U2921 ( .A(n777), .B(n11020), .C(n753), .D(n11262), .Q(n9353) );
  OAI222 U2923 ( .A(n1113), .B(n11018), .C(n1089), .D(n11261), .Q(n9360) );
  OAI222 U2924 ( .A(n1065), .B(n11016), .C(n1041), .D(n11260), .Q(n9359) );
  OAI222 U2925 ( .A(n1017), .B(n11014), .C(n993), .D(n11259), .Q(n9358) );
  OAI222 U2926 ( .A(n969), .B(n11012), .C(n945), .D(n11258), .Q(n9357) );
  OAI222 U2928 ( .A(n1305), .B(n11010), .C(n1281), .D(n11257), .Q(n9364) );
  OAI222 U2929 ( .A(n1257), .B(n11008), .C(n1233), .D(n11256), .Q(n9363) );
  OAI222 U2930 ( .A(n1209), .B(n11006), .C(n1185), .D(n11255), .Q(n9362) );
  OAI222 U2931 ( .A(n1161), .B(n11004), .C(n1137), .D(n11254), .Q(n9361) );
  OAI222 U2933 ( .A(n1497), .B(n11002), .C(n1473), .D(n11253), .Q(n9368) );
  OAI222 U2934 ( .A(n1449), .B(n11000), .C(n1425), .D(n11252), .Q(n9367) );
  OAI222 U2935 ( .A(n1401), .B(n10998), .C(n1377), .D(n11251), .Q(n9366) );
  OAI222 U2936 ( .A(n1353), .B(n10996), .C(n1329), .D(n11250), .Q(n9365) );
  OAI222 U2939 ( .A(n153), .B(n10994), .C(n129), .D(n11249), .Q(n9376) );
  OAI222 U2940 ( .A(n105), .B(n10992), .C(n81), .D(n11248), .Q(n9375) );
  OAI222 U2941 ( .A(n57), .B(n10990), .C(n33), .D(n11247), .Q(n9374) );
  OAI222 U2942 ( .A(n9), .B(n10988), .C(n6129), .D(n11246), .Q(n9373) );
  OAI222 U2944 ( .A(n345), .B(n10986), .C(n321), .D(n11245), .Q(n9380) );
  OAI222 U2945 ( .A(n297), .B(n10984), .C(n273), .D(n11244), .Q(n9379) );
  OAI222 U2946 ( .A(n249), .B(n10982), .C(n225), .D(n11243), .Q(n9378) );
  OAI222 U2947 ( .A(n201), .B(n10980), .C(n177), .D(n11242), .Q(n9377) );
  OAI222 U2949 ( .A(n537), .B(n10978), .C(n513), .D(n11241), .Q(n9384) );
  OAI222 U2950 ( .A(n489), .B(n10976), .C(n465), .D(n11240), .Q(n9383) );
  OAI222 U2951 ( .A(n441), .B(n10974), .C(n417), .D(n11239), .Q(n9382) );
  OAI222 U2952 ( .A(n393), .B(n10972), .C(n369), .D(n11238), .Q(n9381) );
  OAI222 U2954 ( .A(n729), .B(n10970), .C(n705), .D(n11237), .Q(n9388) );
  OAI222 U2955 ( .A(n681), .B(n10968), .C(n657), .D(n11236), .Q(n9387) );
  OAI222 U2956 ( .A(n633), .B(n10966), .C(n609), .D(n11235), .Q(n9386) );
  OAI222 U2957 ( .A(n585), .B(n10964), .C(n561), .D(n11234), .Q(n9385) );
  OAI222 U2961 ( .A(n5529), .B(n10962), .C(n5505), .D(n11233), .Q(n9400) );
  OAI222 U2962 ( .A(n5481), .B(n10960), .C(n5457), .D(n11232), .Q(n9399) );
  OAI222 U2963 ( .A(n5433), .B(n10958), .C(n5409), .D(n11231), .Q(n9398) );
  OAI222 U2964 ( .A(n5385), .B(n10956), .C(n5361), .D(n11230), .Q(n9397) );
  OAI222 U2966 ( .A(n5721), .B(n10954), .C(n5697), .D(n11229), .Q(n9404) );
  OAI222 U2967 ( .A(n5673), .B(n10952), .C(n5649), .D(n11228), .Q(n9403) );
  OAI222 U2968 ( .A(n5625), .B(n10950), .C(n5601), .D(n11227), .Q(n9402) );
  OAI222 U2969 ( .A(n5577), .B(n10948), .C(n5553), .D(n11226), .Q(n9401) );
  OAI222 U2971 ( .A(n5913), .B(n10946), .C(n5889), .D(n11225), .Q(n9408) );
  OAI222 U2972 ( .A(n5865), .B(n10944), .C(n5841), .D(n11224), .Q(n9407) );
  OAI222 U2973 ( .A(n5817), .B(n10942), .C(n5793), .D(n11223), .Q(n9406) );
  OAI222 U2974 ( .A(n5769), .B(n10940), .C(n5745), .D(n11222), .Q(n9405) );
  OAI222 U2976 ( .A(n6105), .B(n10938), .C(n6081), .D(n11221), .Q(n9412) );
  OAI222 U2977 ( .A(n6057), .B(n10936), .C(n6033), .D(n11220), .Q(n9411) );
  OAI222 U2978 ( .A(n6009), .B(n10934), .C(n5985), .D(n11219), .Q(n9410) );
  OAI222 U2979 ( .A(n5961), .B(n10932), .C(n5937), .D(n11218), .Q(n9409) );
  OAI222 U2982 ( .A(n4761), .B(n10930), .C(n4737), .D(n11217), .Q(n9420) );
  OAI222 U2983 ( .A(n4713), .B(n10928), .C(n4689), .D(n11216), .Q(n9419) );
  OAI222 U2984 ( .A(n4665), .B(n10926), .C(n4641), .D(n11215), .Q(n9418) );
  OAI222 U2985 ( .A(n4617), .B(n10924), .C(n4593), .D(n11214), .Q(n9417) );
  OAI222 U2987 ( .A(n4953), .B(n10922), .C(n4929), .D(n11213), .Q(n9424) );
  OAI222 U2988 ( .A(n4905), .B(n10920), .C(n4881), .D(n11212), .Q(n9423) );
  OAI222 U2989 ( .A(n4857), .B(n10918), .C(n4833), .D(n11211), .Q(n9422) );
  OAI222 U2990 ( .A(n4809), .B(n10916), .C(n4785), .D(n11210), .Q(n9421) );
  OAI222 U2992 ( .A(n5145), .B(n10914), .C(n5121), .D(n11209), .Q(n9428) );
  OAI222 U2993 ( .A(n5097), .B(n10912), .C(n5073), .D(n11208), .Q(n9427) );
  OAI222 U2994 ( .A(n5049), .B(n10910), .C(n5025), .D(n11207), .Q(n9426) );
  OAI222 U2995 ( .A(n5001), .B(n10908), .C(n4977), .D(n11206), .Q(n9425) );
  OAI222 U2997 ( .A(n5337), .B(n10906), .C(n5313), .D(n11205), .Q(n9432) );
  OAI222 U2998 ( .A(n5289), .B(n10904), .C(n5265), .D(n11204), .Q(n9431) );
  OAI222 U2999 ( .A(n5241), .B(n10902), .C(n5217), .D(n11203), .Q(n9430) );
  OAI222 U3000 ( .A(n5193), .B(n10900), .C(n5169), .D(n11202), .Q(n9429) );
  OAI222 U3003 ( .A(n3993), .B(n10898), .C(n3969), .D(n11201), .Q(n9440) );
  OAI222 U3004 ( .A(n3945), .B(n10896), .C(n3921), .D(n11200), .Q(n9439) );
  OAI222 U3005 ( .A(n3897), .B(n10894), .C(n3873), .D(n11199), .Q(n9438) );
  OAI222 U3006 ( .A(n3849), .B(n10892), .C(n3825), .D(n11198), .Q(n9437) );
  OAI222 U3008 ( .A(n4185), .B(n10890), .C(n4161), .D(n11197), .Q(n9444) );
  OAI222 U3009 ( .A(n4137), .B(n10888), .C(n4113), .D(n11196), .Q(n9443) );
  OAI222 U3010 ( .A(n4089), .B(n10886), .C(n4065), .D(n11195), .Q(n9442) );
  OAI222 U3011 ( .A(n4041), .B(n10884), .C(n4017), .D(n11194), .Q(n9441) );
  OAI222 U3013 ( .A(n4377), .B(n10882), .C(n4353), .D(n11193), .Q(n9448) );
  OAI222 U3014 ( .A(n4329), .B(n6192), .C(n4305), .D(n11192), .Q(n9447) );
  OAI222 U3015 ( .A(n4281), .B(n6190), .C(n4257), .D(n11191), .Q(n9446) );
  OAI222 U3016 ( .A(n4233), .B(n6188), .C(n4209), .D(n11190), .Q(n9445) );
  OAI222 U3018 ( .A(n4569), .B(n6186), .C(n4545), .D(n11189), .Q(n9452) );
  OAI222 U3019 ( .A(n4521), .B(n6184), .C(n4497), .D(n11188), .Q(n9451) );
  OAI222 U3020 ( .A(n4473), .B(n6182), .C(n4449), .D(n11187), .Q(n9450) );
  OAI222 U3021 ( .A(n4425), .B(n6180), .C(n4401), .D(n11186), .Q(n9449) );
  OAI222 U3024 ( .A(n3225), .B(n6178), .C(n3201), .D(n11185), .Q(n9460) );
  OAI222 U3025 ( .A(n3177), .B(n6176), .C(n3153), .D(n11184), .Q(n9459) );
  OAI222 U3026 ( .A(n3129), .B(n6174), .C(n3105), .D(n11183), .Q(n9458) );
  OAI222 U3027 ( .A(n3081), .B(n6172), .C(n3057), .D(n11182), .Q(n9457) );
  OAI222 U3029 ( .A(n3417), .B(n6170), .C(n3393), .D(n11181), .Q(n9464) );
  OAI222 U3030 ( .A(n3369), .B(n6168), .C(n3345), .D(n11180), .Q(n9463) );
  OAI222 U3031 ( .A(n3321), .B(n6166), .C(n3297), .D(n11179), .Q(n9462) );
  OAI222 U3032 ( .A(n3273), .B(n6164), .C(n3249), .D(n11178), .Q(n9461) );
  OAI222 U3034 ( .A(n3609), .B(n6162), .C(n3585), .D(n11177), .Q(n9468) );
  OAI222 U3035 ( .A(n3561), .B(n6160), .C(n3537), .D(n11176), .Q(n9467) );
  OAI222 U3036 ( .A(n3513), .B(n6158), .C(n3489), .D(n11175), .Q(n9466) );
  OAI222 U3037 ( .A(n3465), .B(n6156), .C(n3441), .D(n11174), .Q(n9465) );
  OAI222 U3039 ( .A(n3801), .B(n6154), .C(n3777), .D(n11173), .Q(n9472) );
  OAI222 U3040 ( .A(n3753), .B(n6152), .C(n3729), .D(n11172), .Q(n9471) );
  OAI222 U3041 ( .A(n3705), .B(n6150), .C(n3681), .D(n11171), .Q(n9470) );
  OAI222 U3042 ( .A(n3657), .B(n6148), .C(n3633), .D(n11170), .Q(n9469) );
  OAI222 U3047 ( .A(n2456), .B(n11090), .C(n2432), .D(n11297), .Q(n9486) );
  OAI222 U3048 ( .A(n2408), .B(n11088), .C(n2384), .D(n11296), .Q(n9485) );
  OAI222 U3049 ( .A(n2360), .B(n11086), .C(n2336), .D(n11295), .Q(n9484) );
  OAI222 U3050 ( .A(n2312), .B(n11084), .C(n2288), .D(n11294), .Q(n9483) );
  OAI222 U3052 ( .A(n2648), .B(n11082), .C(n2624), .D(n11293), .Q(n9490) );
  OAI222 U3053 ( .A(n2600), .B(n11080), .C(n2576), .D(n11292), .Q(n9489) );
  OAI222 U3054 ( .A(n2552), .B(n11078), .C(n2528), .D(n11291), .Q(n9488) );
  OAI222 U3055 ( .A(n2504), .B(n11076), .C(n2480), .D(n11290), .Q(n9487) );
  OAI222 U3057 ( .A(n2840), .B(n11074), .C(n2816), .D(n11289), .Q(n9494) );
  OAI222 U3058 ( .A(n2792), .B(n11072), .C(n2768), .D(n11288), .Q(n9493) );
  OAI222 U3059 ( .A(n2744), .B(n11070), .C(n2720), .D(n11287), .Q(n9492) );
  OAI222 U3060 ( .A(n2696), .B(n11068), .C(n2672), .D(n11286), .Q(n9491) );
  OAI222 U3062 ( .A(n3032), .B(n11066), .C(n3008), .D(n11285), .Q(n9498) );
  OAI222 U3063 ( .A(n2984), .B(n11064), .C(n2960), .D(n11284), .Q(n9497) );
  OAI222 U3064 ( .A(n2936), .B(n11062), .C(n2912), .D(n11283), .Q(n9496) );
  OAI222 U3065 ( .A(n2888), .B(n11060), .C(n2864), .D(n11282), .Q(n9495) );
  OAI222 U3068 ( .A(n1688), .B(n11058), .C(n1664), .D(n11281), .Q(n9506) );
  OAI222 U3069 ( .A(n1640), .B(n11056), .C(n1616), .D(n11280), .Q(n9505) );
  OAI222 U3070 ( .A(n1592), .B(n11054), .C(n1568), .D(n11279), .Q(n9504) );
  OAI222 U3071 ( .A(n1544), .B(n11052), .C(n1520), .D(n11278), .Q(n9503) );
  OAI222 U3073 ( .A(n1880), .B(n11050), .C(n1856), .D(n11277), .Q(n9510) );
  OAI222 U3074 ( .A(n1832), .B(n11048), .C(n1808), .D(n11276), .Q(n9509) );
  OAI222 U3075 ( .A(n1784), .B(n11046), .C(n1760), .D(n11275), .Q(n9508) );
  OAI222 U3076 ( .A(n1736), .B(n11044), .C(n1712), .D(n11274), .Q(n9507) );
  OAI222 U3078 ( .A(n2072), .B(n11042), .C(n2048), .D(n11273), .Q(n9514) );
  OAI222 U3079 ( .A(n2024), .B(n11040), .C(n2000), .D(n11272), .Q(n9513) );
  OAI222 U3080 ( .A(n1976), .B(n11038), .C(n1952), .D(n11271), .Q(n9512) );
  OAI222 U3081 ( .A(n1928), .B(n11036), .C(n1904), .D(n11270), .Q(n9511) );
  OAI222 U3083 ( .A(n2264), .B(n11034), .C(n2240), .D(n11269), .Q(n9518) );
  OAI222 U3084 ( .A(n2216), .B(n11032), .C(n2192), .D(n11268), .Q(n9517) );
  OAI222 U3085 ( .A(n2168), .B(n11030), .C(n2144), .D(n11267), .Q(n9516) );
  OAI222 U3086 ( .A(n2120), .B(n11028), .C(n2096), .D(n11266), .Q(n9515) );
  OAI222 U3089 ( .A(n920), .B(n11026), .C(n896), .D(n11265), .Q(n9526) );
  OAI222 U3090 ( .A(n872), .B(n11024), .C(n848), .D(n11264), .Q(n9525) );
  OAI222 U3091 ( .A(n824), .B(n11022), .C(n800), .D(n11263), .Q(n9524) );
  OAI222 U3092 ( .A(n776), .B(n11020), .C(n752), .D(n11262), .Q(n9523) );
  OAI222 U3094 ( .A(n1112), .B(n11018), .C(n1088), .D(n11261), .Q(n9530) );
  OAI222 U3095 ( .A(n1064), .B(n11016), .C(n1040), .D(n11260), .Q(n9529) );
  OAI222 U3096 ( .A(n1016), .B(n11014), .C(n992), .D(n11259), .Q(n9528) );
  OAI222 U3097 ( .A(n968), .B(n11012), .C(n944), .D(n11258), .Q(n9527) );
  OAI222 U3099 ( .A(n1304), .B(n11010), .C(n1280), .D(n11257), .Q(n9534) );
  OAI222 U3100 ( .A(n1256), .B(n11008), .C(n1232), .D(n11256), .Q(n9533) );
  OAI222 U3101 ( .A(n1208), .B(n11006), .C(n1184), .D(n11255), .Q(n9532) );
  OAI222 U3102 ( .A(n1160), .B(n11004), .C(n1136), .D(n11254), .Q(n9531) );
  OAI222 U3104 ( .A(n1496), .B(n11002), .C(n1472), .D(n11253), .Q(n9538) );
  OAI222 U3105 ( .A(n1448), .B(n11000), .C(n1424), .D(n11252), .Q(n9537) );
  OAI222 U3106 ( .A(n1400), .B(n10998), .C(n1376), .D(n11251), .Q(n9536) );
  OAI222 U3107 ( .A(n1352), .B(n10996), .C(n1328), .D(n11250), .Q(n9535) );
  OAI222 U3110 ( .A(n152), .B(n10994), .C(n128), .D(n11249), .Q(n9546) );
  OAI222 U3111 ( .A(n104), .B(n10992), .C(n80), .D(n11248), .Q(n9545) );
  OAI222 U3112 ( .A(n56), .B(n10990), .C(n32), .D(n11247), .Q(n9544) );
  OAI222 U3113 ( .A(n8), .B(n10988), .C(n6128), .D(n11246), .Q(n9543) );
  OAI222 U3115 ( .A(n344), .B(n10986), .C(n320), .D(n11245), .Q(n9550) );
  OAI222 U3116 ( .A(n296), .B(n10984), .C(n272), .D(n11244), .Q(n9549) );
  OAI222 U3117 ( .A(n248), .B(n10982), .C(n224), .D(n11243), .Q(n9548) );
  OAI222 U3118 ( .A(n200), .B(n10980), .C(n176), .D(n11242), .Q(n9547) );
  OAI222 U3120 ( .A(n536), .B(n10978), .C(n512), .D(n11241), .Q(n9554) );
  OAI222 U3121 ( .A(n488), .B(n10976), .C(n464), .D(n11240), .Q(n9553) );
  OAI222 U3122 ( .A(n440), .B(n10974), .C(n416), .D(n11239), .Q(n9552) );
  OAI222 U3123 ( .A(n392), .B(n10972), .C(n368), .D(n11238), .Q(n9551) );
  OAI222 U3125 ( .A(n728), .B(n10970), .C(n704), .D(n11237), .Q(n9558) );
  OAI222 U3126 ( .A(n680), .B(n10968), .C(n656), .D(n11236), .Q(n9557) );
  OAI222 U3127 ( .A(n632), .B(n10966), .C(n608), .D(n11235), .Q(n9556) );
  OAI222 U3128 ( .A(n584), .B(n10964), .C(n560), .D(n11234), .Q(n9555) );
  OAI222 U3132 ( .A(n5528), .B(n10962), .C(n5504), .D(n11233), .Q(n9570) );
  OAI222 U3133 ( .A(n5480), .B(n10960), .C(n5456), .D(n11232), .Q(n9569) );
  OAI222 U3134 ( .A(n5432), .B(n10958), .C(n5408), .D(n11231), .Q(n9568) );
  OAI222 U3135 ( .A(n5384), .B(n10956), .C(n5360), .D(n11230), .Q(n9567) );
  OAI222 U3137 ( .A(n5720), .B(n10954), .C(n5696), .D(n11229), .Q(n9574) );
  OAI222 U3138 ( .A(n5672), .B(n10952), .C(n5648), .D(n11228), .Q(n9573) );
  OAI222 U3139 ( .A(n5624), .B(n10950), .C(n5600), .D(n11227), .Q(n9572) );
  OAI222 U3140 ( .A(n5576), .B(n10948), .C(n5552), .D(n11226), .Q(n9571) );
  OAI222 U3142 ( .A(n5912), .B(n10946), .C(n5888), .D(n11225), .Q(n9578) );
  OAI222 U3143 ( .A(n5864), .B(n10944), .C(n5840), .D(n11224), .Q(n9577) );
  OAI222 U3144 ( .A(n5816), .B(n10942), .C(n5792), .D(n11223), .Q(n9576) );
  OAI222 U3145 ( .A(n5768), .B(n10940), .C(n5744), .D(n11222), .Q(n9575) );
  OAI222 U3147 ( .A(n6104), .B(n10938), .C(n6080), .D(n11221), .Q(n9582) );
  OAI222 U3148 ( .A(n6056), .B(n10936), .C(n6032), .D(n11220), .Q(n9581) );
  OAI222 U3149 ( .A(n6008), .B(n10934), .C(n5984), .D(n11219), .Q(n9580) );
  OAI222 U3150 ( .A(n5960), .B(n10932), .C(n5936), .D(n11218), .Q(n9579) );
  OAI222 U3153 ( .A(n4760), .B(n10930), .C(n4736), .D(n11217), .Q(n9590) );
  OAI222 U3154 ( .A(n4712), .B(n10928), .C(n4688), .D(n11216), .Q(n9589) );
  OAI222 U3155 ( .A(n4664), .B(n10926), .C(n4640), .D(n11215), .Q(n9588) );
  OAI222 U3156 ( .A(n4616), .B(n10924), .C(n4592), .D(n11214), .Q(n9587) );
  OAI222 U3158 ( .A(n4952), .B(n10922), .C(n4928), .D(n11213), .Q(n9594) );
  OAI222 U3159 ( .A(n4904), .B(n10920), .C(n4880), .D(n11212), .Q(n9593) );
  OAI222 U3160 ( .A(n4856), .B(n10918), .C(n4832), .D(n11211), .Q(n9592) );
  OAI222 U3161 ( .A(n4808), .B(n10916), .C(n4784), .D(n11210), .Q(n9591) );
  OAI222 U3163 ( .A(n5144), .B(n10914), .C(n5120), .D(n11209), .Q(n9598) );
  OAI222 U3164 ( .A(n5096), .B(n10912), .C(n5072), .D(n11208), .Q(n9597) );
  OAI222 U3165 ( .A(n5048), .B(n10910), .C(n5024), .D(n11207), .Q(n9596) );
  OAI222 U3166 ( .A(n5000), .B(n10908), .C(n4976), .D(n11206), .Q(n9595) );
  OAI222 U3168 ( .A(n5336), .B(n10906), .C(n5312), .D(n11205), .Q(n9602) );
  OAI222 U3169 ( .A(n5288), .B(n10904), .C(n5264), .D(n11204), .Q(n9601) );
  OAI222 U3170 ( .A(n5240), .B(n10902), .C(n5216), .D(n11203), .Q(n9600) );
  OAI222 U3171 ( .A(n5192), .B(n10900), .C(n5168), .D(n11202), .Q(n9599) );
  OAI222 U3174 ( .A(n3992), .B(n10898), .C(n3968), .D(n11201), .Q(n9610) );
  OAI222 U3175 ( .A(n3944), .B(n10896), .C(n3920), .D(n11200), .Q(n9609) );
  OAI222 U3176 ( .A(n3896), .B(n10894), .C(n3872), .D(n11199), .Q(n9608) );
  OAI222 U3177 ( .A(n3848), .B(n10892), .C(n3824), .D(n11198), .Q(n9607) );
  OAI222 U3179 ( .A(n4184), .B(n10890), .C(n4160), .D(n11197), .Q(n9614) );
  OAI222 U3180 ( .A(n4136), .B(n10888), .C(n4112), .D(n11196), .Q(n9613) );
  OAI222 U3181 ( .A(n4088), .B(n10886), .C(n4064), .D(n11195), .Q(n9612) );
  OAI222 U3182 ( .A(n4040), .B(n10884), .C(n4016), .D(n11194), .Q(n9611) );
  OAI222 U3184 ( .A(n4376), .B(n10882), .C(n4352), .D(n11193), .Q(n9618) );
  OAI222 U3185 ( .A(n4328), .B(n6192), .C(n4304), .D(n11192), .Q(n9617) );
  OAI222 U3186 ( .A(n4280), .B(n6190), .C(n4256), .D(n11191), .Q(n9616) );
  OAI222 U3187 ( .A(n4232), .B(n6188), .C(n4208), .D(n11190), .Q(n9615) );
  OAI222 U3189 ( .A(n4568), .B(n6186), .C(n4544), .D(n11189), .Q(n9622) );
  OAI222 U3190 ( .A(n4520), .B(n6184), .C(n4496), .D(n11188), .Q(n9621) );
  OAI222 U3191 ( .A(n4472), .B(n6182), .C(n4448), .D(n11187), .Q(n9620) );
  OAI222 U3192 ( .A(n4424), .B(n6180), .C(n4400), .D(n11186), .Q(n9619) );
  OAI222 U3195 ( .A(n3224), .B(n6178), .C(n3200), .D(n11185), .Q(n9630) );
  OAI222 U3196 ( .A(n3176), .B(n6176), .C(n3152), .D(n11184), .Q(n9629) );
  OAI222 U3197 ( .A(n3128), .B(n6174), .C(n3104), .D(n11183), .Q(n9628) );
  OAI222 U3198 ( .A(n3080), .B(n6172), .C(n3056), .D(n11182), .Q(n9627) );
  OAI222 U3200 ( .A(n3416), .B(n6170), .C(n3392), .D(n11181), .Q(n9634) );
  OAI222 U3201 ( .A(n3368), .B(n6168), .C(n3344), .D(n11180), .Q(n9633) );
  OAI222 U3202 ( .A(n3320), .B(n6166), .C(n3296), .D(n11179), .Q(n9632) );
  OAI222 U3203 ( .A(n3272), .B(n6164), .C(n3248), .D(n11178), .Q(n9631) );
  OAI222 U3205 ( .A(n3608), .B(n6162), .C(n3584), .D(n11177), .Q(n9638) );
  OAI222 U3206 ( .A(n3560), .B(n6160), .C(n3536), .D(n11176), .Q(n9637) );
  OAI222 U3207 ( .A(n3512), .B(n6158), .C(n3488), .D(n11175), .Q(n9636) );
  OAI222 U3208 ( .A(n3464), .B(n6156), .C(n3440), .D(n11174), .Q(n9635) );
  OAI222 U3210 ( .A(n3800), .B(n6154), .C(n3776), .D(n11173), .Q(n9642) );
  OAI222 U3211 ( .A(n3752), .B(n6152), .C(n3728), .D(n11172), .Q(n9641) );
  OAI222 U3212 ( .A(n3704), .B(n6150), .C(n3680), .D(n11171), .Q(n9640) );
  OAI222 U3213 ( .A(n3656), .B(n6148), .C(n3632), .D(n11170), .Q(n9639) );
  OAI222 U3218 ( .A(n2455), .B(n11090), .C(n2431), .D(n11297), .Q(n9656) );
  OAI222 U3219 ( .A(n2407), .B(n11088), .C(n2383), .D(n11296), .Q(n9655) );
  OAI222 U3220 ( .A(n2359), .B(n11086), .C(n2335), .D(n11295), .Q(n9654) );
  OAI222 U3221 ( .A(n2311), .B(n11084), .C(n2287), .D(n11294), .Q(n9653) );
  OAI222 U3223 ( .A(n2647), .B(n11082), .C(n2623), .D(n11293), .Q(n9660) );
  OAI222 U3224 ( .A(n2599), .B(n11080), .C(n2575), .D(n11292), .Q(n9659) );
  OAI222 U3225 ( .A(n2551), .B(n11078), .C(n2527), .D(n11291), .Q(n9658) );
  OAI222 U3226 ( .A(n2503), .B(n11076), .C(n2479), .D(n11290), .Q(n9657) );
  OAI222 U3228 ( .A(n2839), .B(n11074), .C(n2815), .D(n11289), .Q(n9664) );
  OAI222 U3229 ( .A(n2791), .B(n11072), .C(n2767), .D(n11288), .Q(n9663) );
  OAI222 U3230 ( .A(n2743), .B(n11070), .C(n2719), .D(n11287), .Q(n9662) );
  OAI222 U3231 ( .A(n2695), .B(n11068), .C(n2671), .D(n11286), .Q(n9661) );
  OAI222 U3233 ( .A(n3031), .B(n11066), .C(n3007), .D(n11285), .Q(n9668) );
  OAI222 U3234 ( .A(n2983), .B(n11064), .C(n2959), .D(n11284), .Q(n9667) );
  OAI222 U3235 ( .A(n2935), .B(n11062), .C(n2911), .D(n11283), .Q(n9666) );
  OAI222 U3236 ( .A(n2887), .B(n11060), .C(n2863), .D(n11282), .Q(n9665) );
  OAI222 U3239 ( .A(n1687), .B(n11058), .C(n1663), .D(n11281), .Q(n9676) );
  OAI222 U3240 ( .A(n1639), .B(n11056), .C(n1615), .D(n11280), .Q(n9675) );
  OAI222 U3241 ( .A(n1591), .B(n11054), .C(n1567), .D(n11279), .Q(n9674) );
  OAI222 U3242 ( .A(n1543), .B(n11052), .C(n1519), .D(n11278), .Q(n9673) );
  OAI222 U3244 ( .A(n1879), .B(n11050), .C(n1855), .D(n11277), .Q(n9680) );
  OAI222 U3245 ( .A(n1831), .B(n11048), .C(n1807), .D(n11276), .Q(n9679) );
  OAI222 U3246 ( .A(n1783), .B(n11046), .C(n1759), .D(n11275), .Q(n9678) );
  OAI222 U3247 ( .A(n1735), .B(n11044), .C(n1711), .D(n11274), .Q(n9677) );
  OAI222 U3249 ( .A(n2071), .B(n11042), .C(n2047), .D(n11273), .Q(n9684) );
  OAI222 U3250 ( .A(n2023), .B(n11040), .C(n1999), .D(n11272), .Q(n9683) );
  OAI222 U3251 ( .A(n1975), .B(n11038), .C(n1951), .D(n11271), .Q(n9682) );
  OAI222 U3252 ( .A(n1927), .B(n11036), .C(n1903), .D(n11270), .Q(n9681) );
  OAI222 U3254 ( .A(n2263), .B(n11034), .C(n2239), .D(n11269), .Q(n9688) );
  OAI222 U3255 ( .A(n2215), .B(n11032), .C(n2191), .D(n11268), .Q(n9687) );
  OAI222 U3256 ( .A(n2167), .B(n11030), .C(n2143), .D(n11267), .Q(n9686) );
  OAI222 U3257 ( .A(n2119), .B(n11028), .C(n2095), .D(n11266), .Q(n9685) );
  OAI222 U3260 ( .A(n919), .B(n11026), .C(n895), .D(n11265), .Q(n9696) );
  OAI222 U3261 ( .A(n871), .B(n11024), .C(n847), .D(n11264), .Q(n9695) );
  OAI222 U3262 ( .A(n823), .B(n11022), .C(n799), .D(n11263), .Q(n9694) );
  OAI222 U3263 ( .A(n775), .B(n11020), .C(n751), .D(n11262), .Q(n9693) );
  OAI222 U3265 ( .A(n1111), .B(n11018), .C(n1087), .D(n11261), .Q(n9700) );
  OAI222 U3266 ( .A(n1063), .B(n11016), .C(n1039), .D(n11260), .Q(n9699) );
  OAI222 U3267 ( .A(n1015), .B(n11014), .C(n991), .D(n11259), .Q(n9698) );
  OAI222 U3268 ( .A(n967), .B(n11012), .C(n943), .D(n11258), .Q(n9697) );
  OAI222 U3270 ( .A(n1303), .B(n11010), .C(n1279), .D(n11257), .Q(n9704) );
  OAI222 U3271 ( .A(n1255), .B(n11008), .C(n1231), .D(n11256), .Q(n9703) );
  OAI222 U3272 ( .A(n1207), .B(n11006), .C(n1183), .D(n11255), .Q(n9702) );
  OAI222 U3273 ( .A(n1159), .B(n11004), .C(n1135), .D(n11254), .Q(n9701) );
  OAI222 U3275 ( .A(n1495), .B(n11002), .C(n1471), .D(n11253), .Q(n9708) );
  OAI222 U3276 ( .A(n1447), .B(n11000), .C(n1423), .D(n11252), .Q(n9707) );
  OAI222 U3277 ( .A(n1399), .B(n10998), .C(n1375), .D(n11251), .Q(n9706) );
  OAI222 U3278 ( .A(n1351), .B(n10996), .C(n1327), .D(n11250), .Q(n9705) );
  OAI222 U3281 ( .A(n151), .B(n10994), .C(n127), .D(n11249), .Q(n9716) );
  OAI222 U3282 ( .A(n103), .B(n10992), .C(n79), .D(n11248), .Q(n9715) );
  OAI222 U3283 ( .A(n55), .B(n10990), .C(n31), .D(n11247), .Q(n9714) );
  OAI222 U3284 ( .A(n7), .B(n10988), .C(n6127), .D(n11246), .Q(n9713) );
  OAI222 U3286 ( .A(n343), .B(n10986), .C(n319), .D(n11245), .Q(n9720) );
  OAI222 U3287 ( .A(n295), .B(n10984), .C(n271), .D(n11244), .Q(n9719) );
  OAI222 U3288 ( .A(n247), .B(n10982), .C(n223), .D(n11243), .Q(n9718) );
  OAI222 U3289 ( .A(n199), .B(n10980), .C(n175), .D(n11242), .Q(n9717) );
  OAI222 U3291 ( .A(n535), .B(n10978), .C(n511), .D(n11241), .Q(n9724) );
  OAI222 U3292 ( .A(n487), .B(n10976), .C(n463), .D(n11240), .Q(n9723) );
  OAI222 U3293 ( .A(n439), .B(n10974), .C(n415), .D(n11239), .Q(n9722) );
  OAI222 U3294 ( .A(n391), .B(n10972), .C(n367), .D(n11238), .Q(n9721) );
  OAI222 U3296 ( .A(n727), .B(n10970), .C(n703), .D(n11237), .Q(n9728) );
  OAI222 U3297 ( .A(n679), .B(n10968), .C(n655), .D(n11236), .Q(n9727) );
  OAI222 U3298 ( .A(n631), .B(n10966), .C(n607), .D(n11235), .Q(n9726) );
  OAI222 U3299 ( .A(n583), .B(n10964), .C(n559), .D(n11234), .Q(n9725) );
  OAI222 U3303 ( .A(n5527), .B(n10962), .C(n5503), .D(n11233), .Q(n9740) );
  OAI222 U3304 ( .A(n5479), .B(n10960), .C(n5455), .D(n11232), .Q(n9739) );
  OAI222 U3305 ( .A(n5431), .B(n10958), .C(n5407), .D(n11231), .Q(n9738) );
  OAI222 U3306 ( .A(n5383), .B(n10956), .C(n5359), .D(n11230), .Q(n9737) );
  OAI222 U3308 ( .A(n5719), .B(n10954), .C(n5695), .D(n11229), .Q(n9744) );
  OAI222 U3309 ( .A(n5671), .B(n10952), .C(n5647), .D(n11228), .Q(n9743) );
  OAI222 U3310 ( .A(n5623), .B(n10950), .C(n5599), .D(n11227), .Q(n9742) );
  OAI222 U3311 ( .A(n5575), .B(n10948), .C(n5551), .D(n11226), .Q(n9741) );
  OAI222 U3313 ( .A(n5911), .B(n10946), .C(n5887), .D(n11225), .Q(n9748) );
  OAI222 U3314 ( .A(n5863), .B(n10944), .C(n5839), .D(n11224), .Q(n9747) );
  OAI222 U3315 ( .A(n5815), .B(n10942), .C(n5791), .D(n11223), .Q(n9746) );
  OAI222 U3316 ( .A(n5767), .B(n10940), .C(n5743), .D(n11222), .Q(n9745) );
  OAI222 U3318 ( .A(n6103), .B(n10938), .C(n6079), .D(n11221), .Q(n9752) );
  OAI222 U3319 ( .A(n6055), .B(n10936), .C(n6031), .D(n11220), .Q(n9751) );
  OAI222 U3320 ( .A(n6007), .B(n10934), .C(n5983), .D(n11219), .Q(n9750) );
  OAI222 U3321 ( .A(n5959), .B(n10932), .C(n5935), .D(n11218), .Q(n9749) );
  OAI222 U3324 ( .A(n4759), .B(n10930), .C(n4735), .D(n11217), .Q(n9760) );
  OAI222 U3325 ( .A(n4711), .B(n10928), .C(n4687), .D(n11216), .Q(n9759) );
  OAI222 U3326 ( .A(n4663), .B(n10926), .C(n4639), .D(n11215), .Q(n9758) );
  OAI222 U3327 ( .A(n4615), .B(n10924), .C(n4591), .D(n11214), .Q(n9757) );
  OAI222 U3329 ( .A(n4951), .B(n10922), .C(n4927), .D(n11213), .Q(n9764) );
  OAI222 U3330 ( .A(n4903), .B(n10920), .C(n4879), .D(n11212), .Q(n9763) );
  OAI222 U3331 ( .A(n4855), .B(n10918), .C(n4831), .D(n11211), .Q(n9762) );
  OAI222 U3332 ( .A(n4807), .B(n10916), .C(n4783), .D(n11210), .Q(n9761) );
  OAI222 U3334 ( .A(n5143), .B(n10914), .C(n5119), .D(n11209), .Q(n9768) );
  OAI222 U3335 ( .A(n5095), .B(n10912), .C(n5071), .D(n11208), .Q(n9767) );
  OAI222 U3336 ( .A(n5047), .B(n10910), .C(n5023), .D(n11207), .Q(n9766) );
  OAI222 U3337 ( .A(n4999), .B(n10908), .C(n4975), .D(n11206), .Q(n9765) );
  OAI222 U3339 ( .A(n5335), .B(n10906), .C(n5311), .D(n11205), .Q(n9772) );
  OAI222 U3340 ( .A(n5287), .B(n10904), .C(n5263), .D(n11204), .Q(n9771) );
  OAI222 U3341 ( .A(n5239), .B(n10902), .C(n5215), .D(n11203), .Q(n9770) );
  OAI222 U3342 ( .A(n5191), .B(n10900), .C(n5167), .D(n11202), .Q(n9769) );
  OAI222 U3345 ( .A(n3991), .B(n10898), .C(n3967), .D(n11201), .Q(n9780) );
  OAI222 U3346 ( .A(n3943), .B(n10896), .C(n3919), .D(n11200), .Q(n9779) );
  OAI222 U3347 ( .A(n3895), .B(n10894), .C(n3871), .D(n11199), .Q(n9778) );
  OAI222 U3348 ( .A(n3847), .B(n10892), .C(n3823), .D(n11198), .Q(n9777) );
  OAI222 U3350 ( .A(n4183), .B(n10890), .C(n4159), .D(n11197), .Q(n9784) );
  OAI222 U3351 ( .A(n4135), .B(n10888), .C(n4111), .D(n11196), .Q(n9783) );
  OAI222 U3352 ( .A(n4087), .B(n10886), .C(n4063), .D(n11195), .Q(n9782) );
  OAI222 U3353 ( .A(n4039), .B(n10884), .C(n4015), .D(n11194), .Q(n9781) );
  OAI222 U3355 ( .A(n4375), .B(n10882), .C(n4351), .D(n11193), .Q(n9788) );
  OAI222 U3356 ( .A(n4327), .B(n6192), .C(n4303), .D(n11192), .Q(n9787) );
  OAI222 U3357 ( .A(n4279), .B(n6190), .C(n4255), .D(n11191), .Q(n9786) );
  OAI222 U3358 ( .A(n4231), .B(n6188), .C(n4207), .D(n11190), .Q(n9785) );
  OAI222 U3360 ( .A(n4567), .B(n6186), .C(n4543), .D(n11189), .Q(n9792) );
  OAI222 U3361 ( .A(n4519), .B(n6184), .C(n4495), .D(n11188), .Q(n9791) );
  OAI222 U3362 ( .A(n4471), .B(n6182), .C(n4447), .D(n11187), .Q(n9790) );
  OAI222 U3363 ( .A(n4423), .B(n6180), .C(n4399), .D(n11186), .Q(n9789) );
  OAI222 U3366 ( .A(n3223), .B(n6178), .C(n3199), .D(n11185), .Q(n9800) );
  OAI222 U3367 ( .A(n3175), .B(n6176), .C(n3151), .D(n11184), .Q(n9799) );
  OAI222 U3368 ( .A(n3127), .B(n6174), .C(n3103), .D(n11183), .Q(n9798) );
  OAI222 U3369 ( .A(n3079), .B(n6172), .C(n3055), .D(n11182), .Q(n9797) );
  OAI222 U3371 ( .A(n3415), .B(n6170), .C(n3391), .D(n11181), .Q(n9804) );
  OAI222 U3372 ( .A(n3367), .B(n6168), .C(n3343), .D(n11180), .Q(n9803) );
  OAI222 U3373 ( .A(n3319), .B(n6166), .C(n3295), .D(n11179), .Q(n9802) );
  OAI222 U3374 ( .A(n3271), .B(n6164), .C(n3247), .D(n11178), .Q(n9801) );
  OAI222 U3376 ( .A(n3607), .B(n6162), .C(n3583), .D(n11177), .Q(n9808) );
  OAI222 U3377 ( .A(n3559), .B(n6160), .C(n3535), .D(n11176), .Q(n9807) );
  OAI222 U3378 ( .A(n3511), .B(n6158), .C(n3487), .D(n11175), .Q(n9806) );
  OAI222 U3379 ( .A(n3463), .B(n6156), .C(n3439), .D(n11174), .Q(n9805) );
  OAI222 U3381 ( .A(n3799), .B(n6154), .C(n3775), .D(n11173), .Q(n9812) );
  OAI222 U3382 ( .A(n3751), .B(n6152), .C(n3727), .D(n11172), .Q(n9811) );
  OAI222 U3383 ( .A(n3703), .B(n6150), .C(n3679), .D(n11171), .Q(n9810) );
  OAI222 U3384 ( .A(n3655), .B(n6148), .C(n3631), .D(n11170), .Q(n9809) );
  OAI222 U3389 ( .A(n2454), .B(n11090), .C(n2430), .D(n11297), .Q(n9826) );
  OAI222 U3390 ( .A(n2406), .B(n11088), .C(n2382), .D(n11296), .Q(n9825) );
  OAI222 U3391 ( .A(n2358), .B(n11086), .C(n2334), .D(n11295), .Q(n9824) );
  OAI222 U3392 ( .A(n2310), .B(n11084), .C(n2286), .D(n11294), .Q(n9823) );
  OAI222 U3394 ( .A(n2646), .B(n11082), .C(n2622), .D(n11293), .Q(n9830) );
  OAI222 U3395 ( .A(n2598), .B(n11080), .C(n2574), .D(n11292), .Q(n9829) );
  OAI222 U3396 ( .A(n2550), .B(n11078), .C(n2526), .D(n11291), .Q(n9828) );
  OAI222 U3397 ( .A(n2502), .B(n11076), .C(n2478), .D(n11290), .Q(n9827) );
  OAI222 U3399 ( .A(n2838), .B(n11074), .C(n2814), .D(n11289), .Q(n9834) );
  OAI222 U3400 ( .A(n2790), .B(n11072), .C(n2766), .D(n11288), .Q(n9833) );
  OAI222 U3401 ( .A(n2742), .B(n11070), .C(n2718), .D(n11287), .Q(n9832) );
  OAI222 U3402 ( .A(n2694), .B(n11068), .C(n2670), .D(n11286), .Q(n9831) );
  OAI222 U3404 ( .A(n3030), .B(n11066), .C(n3006), .D(n11285), .Q(n9838) );
  OAI222 U3405 ( .A(n2982), .B(n11064), .C(n2958), .D(n11284), .Q(n9837) );
  OAI222 U3406 ( .A(n2934), .B(n11062), .C(n2910), .D(n11283), .Q(n9836) );
  OAI222 U3407 ( .A(n2886), .B(n11060), .C(n2862), .D(n11282), .Q(n9835) );
  OAI222 U3410 ( .A(n1686), .B(n11058), .C(n1662), .D(n11281), .Q(n9846) );
  OAI222 U3411 ( .A(n1638), .B(n11056), .C(n1614), .D(n11280), .Q(n9845) );
  OAI222 U3412 ( .A(n1590), .B(n11054), .C(n1566), .D(n11279), .Q(n9844) );
  OAI222 U3413 ( .A(n1542), .B(n11052), .C(n1518), .D(n11278), .Q(n9843) );
  OAI222 U3415 ( .A(n1878), .B(n11050), .C(n1854), .D(n11277), .Q(n9850) );
  OAI222 U3416 ( .A(n1830), .B(n11048), .C(n1806), .D(n11276), .Q(n9849) );
  OAI222 U3417 ( .A(n1782), .B(n11046), .C(n1758), .D(n11275), .Q(n9848) );
  OAI222 U3418 ( .A(n1734), .B(n11044), .C(n1710), .D(n11274), .Q(n9847) );
  OAI222 U3420 ( .A(n2070), .B(n11042), .C(n2046), .D(n11273), .Q(n9854) );
  OAI222 U3421 ( .A(n2022), .B(n11040), .C(n1998), .D(n11272), .Q(n9853) );
  OAI222 U3422 ( .A(n1974), .B(n11038), .C(n1950), .D(n11271), .Q(n9852) );
  OAI222 U3423 ( .A(n1926), .B(n11036), .C(n1902), .D(n11270), .Q(n9851) );
  OAI222 U3425 ( .A(n2262), .B(n11034), .C(n2238), .D(n11269), .Q(n9858) );
  OAI222 U3426 ( .A(n2214), .B(n11032), .C(n2190), .D(n11268), .Q(n9857) );
  OAI222 U3427 ( .A(n2166), .B(n11030), .C(n2142), .D(n11267), .Q(n9856) );
  OAI222 U3428 ( .A(n2118), .B(n11028), .C(n2094), .D(n11266), .Q(n9855) );
  OAI222 U3431 ( .A(n918), .B(n11026), .C(n894), .D(n11265), .Q(n9866) );
  OAI222 U3432 ( .A(n870), .B(n11024), .C(n846), .D(n11264), .Q(n9865) );
  OAI222 U3433 ( .A(n822), .B(n11022), .C(n798), .D(n11263), .Q(n9864) );
  OAI222 U3434 ( .A(n774), .B(n11020), .C(n750), .D(n11262), .Q(n9863) );
  OAI222 U3436 ( .A(n1110), .B(n11018), .C(n1086), .D(n11261), .Q(n9870) );
  OAI222 U3437 ( .A(n1062), .B(n11016), .C(n1038), .D(n11260), .Q(n9869) );
  OAI222 U3438 ( .A(n1014), .B(n11014), .C(n990), .D(n11259), .Q(n9868) );
  OAI222 U3439 ( .A(n966), .B(n11012), .C(n942), .D(n11258), .Q(n9867) );
  OAI222 U3441 ( .A(n1302), .B(n11010), .C(n1278), .D(n11257), .Q(n9874) );
  OAI222 U3442 ( .A(n1254), .B(n11008), .C(n1230), .D(n11256), .Q(n9873) );
  OAI222 U3443 ( .A(n1206), .B(n11006), .C(n1182), .D(n11255), .Q(n9872) );
  OAI222 U3444 ( .A(n1158), .B(n11004), .C(n1134), .D(n11254), .Q(n9871) );
  OAI222 U3446 ( .A(n1494), .B(n11002), .C(n1470), .D(n11253), .Q(n9878) );
  OAI222 U3447 ( .A(n1446), .B(n11000), .C(n1422), .D(n11252), .Q(n9877) );
  OAI222 U3448 ( .A(n1398), .B(n10998), .C(n1374), .D(n11251), .Q(n9876) );
  OAI222 U3449 ( .A(n1350), .B(n10996), .C(n1326), .D(n11250), .Q(n9875) );
  OAI222 U3452 ( .A(n150), .B(n10994), .C(n126), .D(n11249), .Q(n9886) );
  OAI222 U3453 ( .A(n102), .B(n10992), .C(n78), .D(n11248), .Q(n9885) );
  OAI222 U3454 ( .A(n54), .B(n10990), .C(n30), .D(n11247), .Q(n9884) );
  OAI222 U3455 ( .A(n6), .B(n10988), .C(n6126), .D(n11246), .Q(n9883) );
  OAI222 U3457 ( .A(n342), .B(n10986), .C(n318), .D(n11245), .Q(n9890) );
  OAI222 U3458 ( .A(n294), .B(n10984), .C(n270), .D(n11244), .Q(n9889) );
  OAI222 U3459 ( .A(n246), .B(n10982), .C(n222), .D(n11243), .Q(n9888) );
  OAI222 U3460 ( .A(n198), .B(n10980), .C(n174), .D(n11242), .Q(n9887) );
  OAI222 U3462 ( .A(n534), .B(n10978), .C(n510), .D(n11241), .Q(n9894) );
  OAI222 U3463 ( .A(n486), .B(n10976), .C(n462), .D(n11240), .Q(n9893) );
  OAI222 U3464 ( .A(n438), .B(n10974), .C(n414), .D(n11239), .Q(n9892) );
  OAI222 U3465 ( .A(n390), .B(n10972), .C(n366), .D(n11238), .Q(n9891) );
  OAI222 U3467 ( .A(n726), .B(n10970), .C(n702), .D(n11237), .Q(n9898) );
  OAI222 U3468 ( .A(n678), .B(n10968), .C(n654), .D(n11236), .Q(n9897) );
  OAI222 U3469 ( .A(n630), .B(n10966), .C(n606), .D(n11235), .Q(n9896) );
  OAI222 U3470 ( .A(n582), .B(n10964), .C(n558), .D(n11234), .Q(n9895) );
  OAI222 U3474 ( .A(n5526), .B(n10962), .C(n5502), .D(n11233), .Q(n9910) );
  OAI222 U3475 ( .A(n5478), .B(n10960), .C(n5454), .D(n11232), .Q(n9909) );
  OAI222 U3476 ( .A(n5430), .B(n10958), .C(n5406), .D(n11231), .Q(n9908) );
  OAI222 U3477 ( .A(n5382), .B(n10956), .C(n5358), .D(n11230), .Q(n9907) );
  OAI222 U3479 ( .A(n5718), .B(n10954), .C(n5694), .D(n11229), .Q(n9914) );
  OAI222 U3480 ( .A(n5670), .B(n10952), .C(n5646), .D(n11228), .Q(n9913) );
  OAI222 U3481 ( .A(n5622), .B(n10950), .C(n5598), .D(n11227), .Q(n9912) );
  OAI222 U3482 ( .A(n5574), .B(n10948), .C(n5550), .D(n11226), .Q(n9911) );
  OAI222 U3484 ( .A(n5910), .B(n10946), .C(n5886), .D(n11225), .Q(n9918) );
  OAI222 U3485 ( .A(n5862), .B(n10944), .C(n5838), .D(n11224), .Q(n9917) );
  OAI222 U3486 ( .A(n5814), .B(n10942), .C(n5790), .D(n11223), .Q(n9916) );
  OAI222 U3487 ( .A(n5766), .B(n10940), .C(n5742), .D(n11222), .Q(n9915) );
  OAI222 U3489 ( .A(n6102), .B(n10938), .C(n6078), .D(n11221), .Q(n9922) );
  OAI222 U3490 ( .A(n6054), .B(n10936), .C(n6030), .D(n11220), .Q(n9921) );
  OAI222 U3491 ( .A(n6006), .B(n10934), .C(n5982), .D(n11219), .Q(n9920) );
  OAI222 U3492 ( .A(n5958), .B(n10932), .C(n5934), .D(n11218), .Q(n9919) );
  OAI222 U3495 ( .A(n4758), .B(n10930), .C(n4734), .D(n11217), .Q(n9930) );
  OAI222 U3496 ( .A(n4710), .B(n10928), .C(n4686), .D(n11216), .Q(n9929) );
  OAI222 U3497 ( .A(n4662), .B(n10926), .C(n4638), .D(n11215), .Q(n9928) );
  OAI222 U3498 ( .A(n4614), .B(n10924), .C(n4590), .D(n11214), .Q(n9927) );
  OAI222 U3500 ( .A(n4950), .B(n10922), .C(n4926), .D(n11213), .Q(n9934) );
  OAI222 U3501 ( .A(n4902), .B(n10920), .C(n4878), .D(n11212), .Q(n9933) );
  OAI222 U3502 ( .A(n4854), .B(n10918), .C(n4830), .D(n11211), .Q(n9932) );
  OAI222 U3503 ( .A(n4806), .B(n10916), .C(n4782), .D(n11210), .Q(n9931) );
  OAI222 U3505 ( .A(n5142), .B(n10914), .C(n5118), .D(n11209), .Q(n9938) );
  OAI222 U3506 ( .A(n5094), .B(n10912), .C(n5070), .D(n11208), .Q(n9937) );
  OAI222 U3507 ( .A(n5046), .B(n10910), .C(n5022), .D(n11207), .Q(n9936) );
  OAI222 U3508 ( .A(n4998), .B(n10908), .C(n4974), .D(n11206), .Q(n9935) );
  OAI222 U3510 ( .A(n5334), .B(n10906), .C(n5310), .D(n11205), .Q(n9942) );
  OAI222 U3511 ( .A(n5286), .B(n10904), .C(n5262), .D(n11204), .Q(n9941) );
  OAI222 U3512 ( .A(n5238), .B(n10902), .C(n5214), .D(n11203), .Q(n9940) );
  OAI222 U3513 ( .A(n5190), .B(n10900), .C(n5166), .D(n11202), .Q(n9939) );
  OAI222 U3516 ( .A(n3990), .B(n10898), .C(n3966), .D(n11201), .Q(n9950) );
  OAI222 U3517 ( .A(n3942), .B(n10896), .C(n3918), .D(n11200), .Q(n9949) );
  OAI222 U3518 ( .A(n3894), .B(n10894), .C(n3870), .D(n11199), .Q(n9948) );
  OAI222 U3519 ( .A(n3846), .B(n10892), .C(n3822), .D(n11198), .Q(n9947) );
  OAI222 U3521 ( .A(n4182), .B(n10890), .C(n4158), .D(n11197), .Q(n9954) );
  OAI222 U3522 ( .A(n4134), .B(n10888), .C(n4110), .D(n11196), .Q(n9953) );
  OAI222 U3523 ( .A(n4086), .B(n10886), .C(n4062), .D(n11195), .Q(n9952) );
  OAI222 U3524 ( .A(n4038), .B(n10884), .C(n4014), .D(n11194), .Q(n9951) );
  OAI222 U3526 ( .A(n4374), .B(n10882), .C(n4350), .D(n11193), .Q(n9958) );
  OAI222 U3527 ( .A(n4326), .B(n6192), .C(n4302), .D(n11192), .Q(n9957) );
  OAI222 U3528 ( .A(n4278), .B(n6190), .C(n4254), .D(n11191), .Q(n9956) );
  OAI222 U3529 ( .A(n4230), .B(n6188), .C(n4206), .D(n11190), .Q(n9955) );
  OAI222 U3531 ( .A(n4566), .B(n6186), .C(n4542), .D(n11189), .Q(n9962) );
  OAI222 U3532 ( .A(n4518), .B(n6184), .C(n4494), .D(n11188), .Q(n9961) );
  OAI222 U3533 ( .A(n4470), .B(n6182), .C(n4446), .D(n11187), .Q(n9960) );
  OAI222 U3534 ( .A(n4422), .B(n6180), .C(n4398), .D(n11186), .Q(n9959) );
  OAI222 U3537 ( .A(n3222), .B(n6178), .C(n3198), .D(n11185), .Q(n9970) );
  OAI222 U3538 ( .A(n3174), .B(n6176), .C(n3150), .D(n11184), .Q(n9969) );
  OAI222 U3539 ( .A(n3126), .B(n6174), .C(n3102), .D(n11183), .Q(n9968) );
  OAI222 U3540 ( .A(n3078), .B(n6172), .C(n3054), .D(n11182), .Q(n9967) );
  OAI222 U3542 ( .A(n3414), .B(n6170), .C(n3390), .D(n11181), .Q(n9974) );
  OAI222 U3543 ( .A(n3366), .B(n6168), .C(n3342), .D(n11180), .Q(n9973) );
  OAI222 U3544 ( .A(n3318), .B(n6166), .C(n3294), .D(n11179), .Q(n9972) );
  OAI222 U3545 ( .A(n3270), .B(n6164), .C(n3246), .D(n11178), .Q(n9971) );
  OAI222 U3547 ( .A(n3606), .B(n6162), .C(n3582), .D(n11177), .Q(n9978) );
  OAI222 U3548 ( .A(n3558), .B(n6160), .C(n3534), .D(n11176), .Q(n9977) );
  OAI222 U3549 ( .A(n3510), .B(n6158), .C(n3486), .D(n11175), .Q(n9976) );
  OAI222 U3550 ( .A(n3462), .B(n6156), .C(n3438), .D(n11174), .Q(n9975) );
  OAI222 U3552 ( .A(n3798), .B(n6154), .C(n3774), .D(n11173), .Q(n9982) );
  OAI222 U3553 ( .A(n3750), .B(n6152), .C(n3726), .D(n11172), .Q(n9981) );
  OAI222 U3554 ( .A(n3702), .B(n6150), .C(n3678), .D(n11171), .Q(n9980) );
  OAI222 U3555 ( .A(n3654), .B(n6148), .C(n3630), .D(n11170), .Q(n9979) );
  OAI222 U3560 ( .A(n2453), .B(n11090), .C(n2429), .D(n11297), .Q(n9996) );
  OAI222 U3561 ( .A(n2405), .B(n11088), .C(n2381), .D(n11296), .Q(n9995) );
  OAI222 U3562 ( .A(n2357), .B(n11086), .C(n2333), .D(n11295), .Q(n9994) );
  OAI222 U3563 ( .A(n2309), .B(n11084), .C(n2285), .D(n11294), .Q(n9993) );
  OAI222 U3565 ( .A(n2645), .B(n11082), .C(n2621), .D(n11293), .Q(n10000) );
  OAI222 U3566 ( .A(n2597), .B(n11080), .C(n2573), .D(n11292), .Q(n9999) );
  OAI222 U3567 ( .A(n2549), .B(n11078), .C(n2525), .D(n11291), .Q(n9998) );
  OAI222 U3568 ( .A(n2501), .B(n11076), .C(n2477), .D(n11290), .Q(n9997) );
  OAI222 U3570 ( .A(n2837), .B(n11074), .C(n2813), .D(n11289), .Q(n10004) );
  OAI222 U3571 ( .A(n2789), .B(n11072), .C(n2765), .D(n11288), .Q(n10003) );
  OAI222 U3572 ( .A(n2741), .B(n11070), .C(n2717), .D(n11287), .Q(n10002) );
  OAI222 U3573 ( .A(n2693), .B(n11068), .C(n2669), .D(n11286), .Q(n10001) );
  OAI222 U3575 ( .A(n3029), .B(n11066), .C(n3005), .D(n11285), .Q(n10008) );
  OAI222 U3576 ( .A(n2981), .B(n11064), .C(n2957), .D(n11284), .Q(n10007) );
  OAI222 U3577 ( .A(n2933), .B(n11062), .C(n2909), .D(n11283), .Q(n10006) );
  OAI222 U3578 ( .A(n2885), .B(n11060), .C(n2861), .D(n11282), .Q(n10005) );
  OAI222 U3581 ( .A(n1685), .B(n11058), .C(n1661), .D(n11281), .Q(n10016) );
  OAI222 U3582 ( .A(n1637), .B(n11056), .C(n1613), .D(n11280), .Q(n10015) );
  OAI222 U3583 ( .A(n1589), .B(n11054), .C(n1565), .D(n11279), .Q(n10014) );
  OAI222 U3584 ( .A(n1541), .B(n11052), .C(n1517), .D(n11278), .Q(n10013) );
  OAI222 U3586 ( .A(n1877), .B(n11050), .C(n1853), .D(n11277), .Q(n10020) );
  OAI222 U3587 ( .A(n1829), .B(n11048), .C(n1805), .D(n11276), .Q(n10019) );
  OAI222 U3588 ( .A(n1781), .B(n11046), .C(n1757), .D(n11275), .Q(n10018) );
  OAI222 U3589 ( .A(n1733), .B(n11044), .C(n1709), .D(n11274), .Q(n10017) );
  OAI222 U3591 ( .A(n2069), .B(n11042), .C(n2045), .D(n11273), .Q(n10024) );
  OAI222 U3592 ( .A(n2021), .B(n11040), .C(n1997), .D(n11272), .Q(n10023) );
  OAI222 U3593 ( .A(n1973), .B(n11038), .C(n1949), .D(n11271), .Q(n10022) );
  OAI222 U3594 ( .A(n1925), .B(n11036), .C(n1901), .D(n11270), .Q(n10021) );
  OAI222 U3596 ( .A(n2261), .B(n11034), .C(n2237), .D(n11269), .Q(n10028) );
  OAI222 U3597 ( .A(n2213), .B(n11032), .C(n2189), .D(n11268), .Q(n10027) );
  OAI222 U3598 ( .A(n2165), .B(n11030), .C(n2141), .D(n11267), .Q(n10026) );
  OAI222 U3599 ( .A(n2117), .B(n11028), .C(n2093), .D(n11266), .Q(n10025) );
  OAI222 U3602 ( .A(n917), .B(n11026), .C(n893), .D(n11265), .Q(n10036) );
  OAI222 U3603 ( .A(n869), .B(n11024), .C(n845), .D(n11264), .Q(n10035) );
  OAI222 U3604 ( .A(n821), .B(n11022), .C(n797), .D(n11263), .Q(n10034) );
  OAI222 U3605 ( .A(n773), .B(n11020), .C(n749), .D(n11262), .Q(n10033) );
  OAI222 U3607 ( .A(n1109), .B(n11018), .C(n1085), .D(n11261), .Q(n10040) );
  OAI222 U3608 ( .A(n1061), .B(n11016), .C(n1037), .D(n11260), .Q(n10039) );
  OAI222 U3609 ( .A(n1013), .B(n11014), .C(n989), .D(n11259), .Q(n10038) );
  OAI222 U3610 ( .A(n965), .B(n11012), .C(n941), .D(n11258), .Q(n10037) );
  OAI222 U3612 ( .A(n1301), .B(n11010), .C(n1277), .D(n11257), .Q(n10044) );
  OAI222 U3613 ( .A(n1253), .B(n11008), .C(n1229), .D(n11256), .Q(n10043) );
  OAI222 U3614 ( .A(n1205), .B(n11006), .C(n1181), .D(n11255), .Q(n10042) );
  OAI222 U3615 ( .A(n1157), .B(n11004), .C(n1133), .D(n11254), .Q(n10041) );
  OAI222 U3617 ( .A(n1493), .B(n11002), .C(n1469), .D(n11253), .Q(n10048) );
  OAI222 U3618 ( .A(n1445), .B(n11000), .C(n1421), .D(n11252), .Q(n10047) );
  OAI222 U3619 ( .A(n1397), .B(n10998), .C(n1373), .D(n11251), .Q(n10046) );
  OAI222 U3620 ( .A(n1349), .B(n10996), .C(n1325), .D(n11250), .Q(n10045) );
  OAI222 U3623 ( .A(n149), .B(n10994), .C(n125), .D(n11249), .Q(n10056) );
  OAI222 U3624 ( .A(n101), .B(n10992), .C(n77), .D(n11248), .Q(n10055) );
  OAI222 U3625 ( .A(n53), .B(n10990), .C(n29), .D(n11247), .Q(n10054) );
  OAI222 U3626 ( .A(n5), .B(n10988), .C(n6125), .D(n11246), .Q(n10053) );
  OAI222 U3628 ( .A(n341), .B(n10986), .C(n317), .D(n11245), .Q(n10060) );
  OAI222 U3629 ( .A(n293), .B(n10984), .C(n269), .D(n11244), .Q(n10059) );
  OAI222 U3630 ( .A(n245), .B(n10982), .C(n221), .D(n11243), .Q(n10058) );
  OAI222 U3631 ( .A(n197), .B(n10980), .C(n173), .D(n11242), .Q(n10057) );
  OAI222 U3633 ( .A(n533), .B(n10978), .C(n509), .D(n11241), .Q(n10064) );
  OAI222 U3634 ( .A(n485), .B(n10976), .C(n461), .D(n11240), .Q(n10063) );
  OAI222 U3635 ( .A(n437), .B(n10974), .C(n413), .D(n11239), .Q(n10062) );
  OAI222 U3636 ( .A(n389), .B(n10972), .C(n365), .D(n11238), .Q(n10061) );
  OAI222 U3638 ( .A(n725), .B(n10970), .C(n701), .D(n11237), .Q(n10068) );
  OAI222 U3639 ( .A(n677), .B(n10968), .C(n653), .D(n11236), .Q(n10067) );
  OAI222 U3640 ( .A(n629), .B(n10966), .C(n605), .D(n11235), .Q(n10066) );
  OAI222 U3641 ( .A(n581), .B(n10964), .C(n557), .D(n11234), .Q(n10065) );
  OAI222 U3645 ( .A(n5525), .B(n10962), .C(n5501), .D(n11233), .Q(n10080) );
  OAI222 U3646 ( .A(n5477), .B(n10960), .C(n5453), .D(n11232), .Q(n10079) );
  OAI222 U3647 ( .A(n5429), .B(n10958), .C(n5405), .D(n11231), .Q(n10078) );
  OAI222 U3648 ( .A(n5381), .B(n10956), .C(n5357), .D(n11230), .Q(n10077) );
  OAI222 U3650 ( .A(n5717), .B(n10954), .C(n5693), .D(n11229), .Q(n10084) );
  OAI222 U3651 ( .A(n5669), .B(n10952), .C(n5645), .D(n11228), .Q(n10083) );
  OAI222 U3652 ( .A(n5621), .B(n10950), .C(n5597), .D(n11227), .Q(n10082) );
  OAI222 U3653 ( .A(n5573), .B(n10948), .C(n5549), .D(n11226), .Q(n10081) );
  OAI222 U3655 ( .A(n5909), .B(n10946), .C(n5885), .D(n11225), .Q(n10088) );
  OAI222 U3656 ( .A(n5861), .B(n10944), .C(n5837), .D(n11224), .Q(n10087) );
  OAI222 U3657 ( .A(n5813), .B(n10942), .C(n5789), .D(n11223), .Q(n10086) );
  OAI222 U3658 ( .A(n5765), .B(n10940), .C(n5741), .D(n11222), .Q(n10085) );
  OAI222 U3660 ( .A(n6101), .B(n10938), .C(n6077), .D(n11221), .Q(n10092) );
  OAI222 U3661 ( .A(n6053), .B(n10936), .C(n6029), .D(n11220), .Q(n10091) );
  OAI222 U3662 ( .A(n6005), .B(n10934), .C(n5981), .D(n11219), .Q(n10090) );
  OAI222 U3663 ( .A(n5957), .B(n10932), .C(n5933), .D(n11218), .Q(n10089) );
  OAI222 U3666 ( .A(n4757), .B(n10930), .C(n4733), .D(n11217), .Q(n10100) );
  OAI222 U3667 ( .A(n4709), .B(n10928), .C(n4685), .D(n11216), .Q(n10099) );
  OAI222 U3668 ( .A(n4661), .B(n10926), .C(n4637), .D(n11215), .Q(n10098) );
  OAI222 U3669 ( .A(n4613), .B(n10924), .C(n4589), .D(n11214), .Q(n10097) );
  OAI222 U3671 ( .A(n4949), .B(n10922), .C(n4925), .D(n11213), .Q(n10104) );
  OAI222 U3672 ( .A(n4901), .B(n10920), .C(n4877), .D(n11212), .Q(n10103) );
  OAI222 U3673 ( .A(n4853), .B(n10918), .C(n4829), .D(n11211), .Q(n10102) );
  OAI222 U3674 ( .A(n4805), .B(n10916), .C(n4781), .D(n11210), .Q(n10101) );
  OAI222 U3676 ( .A(n5141), .B(n10914), .C(n5117), .D(n11209), .Q(n10108) );
  OAI222 U3677 ( .A(n5093), .B(n10912), .C(n5069), .D(n11208), .Q(n10107) );
  OAI222 U3678 ( .A(n5045), .B(n10910), .C(n5021), .D(n11207), .Q(n10106) );
  OAI222 U3679 ( .A(n4997), .B(n10908), .C(n4973), .D(n11206), .Q(n10105) );
  OAI222 U3681 ( .A(n5333), .B(n10906), .C(n5309), .D(n11205), .Q(n10112) );
  OAI222 U3682 ( .A(n5285), .B(n10904), .C(n5261), .D(n11204), .Q(n10111) );
  OAI222 U3683 ( .A(n5237), .B(n10902), .C(n5213), .D(n11203), .Q(n10110) );
  OAI222 U3684 ( .A(n5189), .B(n10900), .C(n5165), .D(n11202), .Q(n10109) );
  OAI222 U3687 ( .A(n3989), .B(n10898), .C(n3965), .D(n11201), .Q(n10120) );
  OAI222 U3688 ( .A(n3941), .B(n10896), .C(n3917), .D(n11200), .Q(n10119) );
  OAI222 U3689 ( .A(n3893), .B(n10894), .C(n3869), .D(n11199), .Q(n10118) );
  OAI222 U3690 ( .A(n3845), .B(n10892), .C(n3821), .D(n11198), .Q(n10117) );
  OAI222 U3692 ( .A(n4181), .B(n10890), .C(n4157), .D(n11197), .Q(n10124) );
  OAI222 U3693 ( .A(n4133), .B(n10888), .C(n4109), .D(n11196), .Q(n10123) );
  OAI222 U3694 ( .A(n4085), .B(n10886), .C(n4061), .D(n11195), .Q(n10122) );
  OAI222 U3695 ( .A(n4037), .B(n10884), .C(n4013), .D(n11194), .Q(n10121) );
  OAI222 U3697 ( .A(n4373), .B(n10882), .C(n4349), .D(n11193), .Q(n10128) );
  OAI222 U3698 ( .A(n4325), .B(n6192), .C(n4301), .D(n11192), .Q(n10127) );
  OAI222 U3699 ( .A(n4277), .B(n6190), .C(n4253), .D(n11191), .Q(n10126) );
  OAI222 U3700 ( .A(n4229), .B(n6188), .C(n4205), .D(n11190), .Q(n10125) );
  OAI222 U3702 ( .A(n4565), .B(n6186), .C(n4541), .D(n11189), .Q(n10132) );
  OAI222 U3703 ( .A(n4517), .B(n6184), .C(n4493), .D(n11188), .Q(n10131) );
  OAI222 U3704 ( .A(n4469), .B(n6182), .C(n4445), .D(n11187), .Q(n10130) );
  OAI222 U3705 ( .A(n4421), .B(n6180), .C(n4397), .D(n11186), .Q(n10129) );
  OAI222 U3708 ( .A(n3221), .B(n6178), .C(n3197), .D(n11185), .Q(n10140) );
  OAI222 U3709 ( .A(n3173), .B(n6176), .C(n3149), .D(n11184), .Q(n10139) );
  OAI222 U3710 ( .A(n3125), .B(n6174), .C(n3101), .D(n11183), .Q(n10138) );
  OAI222 U3711 ( .A(n3077), .B(n6172), .C(n3053), .D(n11182), .Q(n10137) );
  OAI222 U3713 ( .A(n3413), .B(n6170), .C(n3389), .D(n11181), .Q(n10144) );
  OAI222 U3714 ( .A(n3365), .B(n6168), .C(n3341), .D(n11180), .Q(n10143) );
  OAI222 U3715 ( .A(n3317), .B(n6166), .C(n3293), .D(n11179), .Q(n10142) );
  OAI222 U3716 ( .A(n3269), .B(n6164), .C(n3245), .D(n11178), .Q(n10141) );
  OAI222 U3718 ( .A(n3605), .B(n6162), .C(n3581), .D(n11177), .Q(n10148) );
  OAI222 U3719 ( .A(n3557), .B(n6160), .C(n3533), .D(n11176), .Q(n10147) );
  OAI222 U3720 ( .A(n3509), .B(n6158), .C(n3485), .D(n11175), .Q(n10146) );
  OAI222 U3721 ( .A(n3461), .B(n6156), .C(n3437), .D(n11174), .Q(n10145) );
  OAI222 U3723 ( .A(n3797), .B(n6154), .C(n3773), .D(n11173), .Q(n10152) );
  OAI222 U3724 ( .A(n3749), .B(n6152), .C(n3725), .D(n11172), .Q(n10151) );
  OAI222 U3725 ( .A(n3701), .B(n6150), .C(n3677), .D(n11171), .Q(n10150) );
  OAI222 U3726 ( .A(n3653), .B(n6148), .C(n3629), .D(n11170), .Q(n10149) );
  OAI222 U3731 ( .A(n2452), .B(n11090), .C(n2428), .D(n11297), .Q(n10166) );
  OAI222 U3732 ( .A(n2404), .B(n11088), .C(n2380), .D(n11296), .Q(n10165) );
  OAI222 U3733 ( .A(n2356), .B(n11086), .C(n2332), .D(n11295), .Q(n10164) );
  OAI222 U3734 ( .A(n2308), .B(n11084), .C(n2284), .D(n11294), .Q(n10163) );
  OAI222 U3736 ( .A(n2644), .B(n11082), .C(n2620), .D(n11293), .Q(n10170) );
  OAI222 U3737 ( .A(n2596), .B(n11080), .C(n2572), .D(n11292), .Q(n10169) );
  OAI222 U3738 ( .A(n2548), .B(n11078), .C(n2524), .D(n11291), .Q(n10168) );
  OAI222 U3739 ( .A(n2500), .B(n11076), .C(n2476), .D(n11290), .Q(n10167) );
  OAI222 U3741 ( .A(n2836), .B(n11074), .C(n2812), .D(n11289), .Q(n10174) );
  OAI222 U3742 ( .A(n2788), .B(n11072), .C(n2764), .D(n11288), .Q(n10173) );
  OAI222 U3743 ( .A(n2740), .B(n11070), .C(n2716), .D(n11287), .Q(n10172) );
  OAI222 U3744 ( .A(n2692), .B(n11068), .C(n2668), .D(n11286), .Q(n10171) );
  OAI222 U3746 ( .A(n3028), .B(n11066), .C(n3004), .D(n11285), .Q(n10178) );
  OAI222 U3747 ( .A(n2980), .B(n11064), .C(n2956), .D(n11284), .Q(n10177) );
  OAI222 U3748 ( .A(n2932), .B(n11062), .C(n2908), .D(n11283), .Q(n10176) );
  OAI222 U3749 ( .A(n2884), .B(n11060), .C(n2860), .D(n11282), .Q(n10175) );
  OAI222 U3752 ( .A(n1684), .B(n11058), .C(n1660), .D(n11281), .Q(n10186) );
  OAI222 U3753 ( .A(n1636), .B(n11056), .C(n1612), .D(n11280), .Q(n10185) );
  OAI222 U3754 ( .A(n1588), .B(n11054), .C(n1564), .D(n11279), .Q(n10184) );
  OAI222 U3755 ( .A(n1540), .B(n11052), .C(n1516), .D(n11278), .Q(n10183) );
  OAI222 U3757 ( .A(n1876), .B(n11050), .C(n1852), .D(n11277), .Q(n10190) );
  OAI222 U3758 ( .A(n1828), .B(n11048), .C(n1804), .D(n11276), .Q(n10189) );
  OAI222 U3759 ( .A(n1780), .B(n11046), .C(n1756), .D(n11275), .Q(n10188) );
  OAI222 U3760 ( .A(n1732), .B(n11044), .C(n1708), .D(n11274), .Q(n10187) );
  OAI222 U3762 ( .A(n2068), .B(n11042), .C(n2044), .D(n11273), .Q(n10194) );
  OAI222 U3763 ( .A(n2020), .B(n11040), .C(n1996), .D(n11272), .Q(n10193) );
  OAI222 U3764 ( .A(n1972), .B(n11038), .C(n1948), .D(n11271), .Q(n10192) );
  OAI222 U3765 ( .A(n1924), .B(n11036), .C(n1900), .D(n11270), .Q(n10191) );
  OAI222 U3767 ( .A(n2260), .B(n11034), .C(n2236), .D(n11269), .Q(n10198) );
  OAI222 U3768 ( .A(n2212), .B(n11032), .C(n2188), .D(n11268), .Q(n10197) );
  OAI222 U3769 ( .A(n2164), .B(n11030), .C(n2140), .D(n11267), .Q(n10196) );
  OAI222 U3770 ( .A(n2116), .B(n11028), .C(n2092), .D(n11266), .Q(n10195) );
  OAI222 U3773 ( .A(n916), .B(n11026), .C(n892), .D(n11265), .Q(n10206) );
  OAI222 U3774 ( .A(n868), .B(n11024), .C(n844), .D(n11264), .Q(n10205) );
  OAI222 U3775 ( .A(n820), .B(n11022), .C(n796), .D(n11263), .Q(n10204) );
  OAI222 U3776 ( .A(n772), .B(n11020), .C(n748), .D(n11262), .Q(n10203) );
  OAI222 U3778 ( .A(n1108), .B(n11018), .C(n1084), .D(n11261), .Q(n10210) );
  OAI222 U3779 ( .A(n1060), .B(n11016), .C(n1036), .D(n11260), .Q(n10209) );
  OAI222 U3780 ( .A(n1012), .B(n11014), .C(n988), .D(n11259), .Q(n10208) );
  OAI222 U3781 ( .A(n964), .B(n11012), .C(n940), .D(n11258), .Q(n10207) );
  OAI222 U3783 ( .A(n1300), .B(n11010), .C(n1276), .D(n11257), .Q(n10214) );
  OAI222 U3784 ( .A(n1252), .B(n11008), .C(n1228), .D(n11256), .Q(n10213) );
  OAI222 U3785 ( .A(n1204), .B(n11006), .C(n1180), .D(n11255), .Q(n10212) );
  OAI222 U3786 ( .A(n1156), .B(n11004), .C(n1132), .D(n11254), .Q(n10211) );
  OAI222 U3788 ( .A(n1492), .B(n11002), .C(n1468), .D(n11253), .Q(n10218) );
  OAI222 U3789 ( .A(n1444), .B(n11000), .C(n1420), .D(n11252), .Q(n10217) );
  OAI222 U3790 ( .A(n1396), .B(n10998), .C(n1372), .D(n11251), .Q(n10216) );
  OAI222 U3791 ( .A(n1348), .B(n10996), .C(n1324), .D(n11250), .Q(n10215) );
  OAI222 U3794 ( .A(n148), .B(n10994), .C(n124), .D(n11249), .Q(n10226) );
  OAI222 U3795 ( .A(n100), .B(n10992), .C(n76), .D(n11248), .Q(n10225) );
  OAI222 U3796 ( .A(n52), .B(n10990), .C(n28), .D(n11247), .Q(n10224) );
  OAI222 U3797 ( .A(n4), .B(n10988), .C(n6124), .D(n11246), .Q(n10223) );
  OAI222 U3799 ( .A(n340), .B(n10986), .C(n316), .D(n11245), .Q(n10230) );
  OAI222 U3800 ( .A(n292), .B(n10984), .C(n268), .D(n11244), .Q(n10229) );
  OAI222 U3801 ( .A(n244), .B(n10982), .C(n220), .D(n11243), .Q(n10228) );
  OAI222 U3802 ( .A(n196), .B(n10980), .C(n172), .D(n11242), .Q(n10227) );
  OAI222 U3804 ( .A(n532), .B(n10978), .C(n508), .D(n11241), .Q(n10234) );
  OAI222 U3805 ( .A(n484), .B(n10976), .C(n460), .D(n11240), .Q(n10233) );
  OAI222 U3806 ( .A(n436), .B(n10974), .C(n412), .D(n11239), .Q(n10232) );
  OAI222 U3807 ( .A(n388), .B(n10972), .C(n364), .D(n11238), .Q(n10231) );
  OAI222 U3809 ( .A(n724), .B(n10970), .C(n700), .D(n11237), .Q(n10238) );
  OAI222 U3810 ( .A(n676), .B(n10968), .C(n652), .D(n11236), .Q(n10237) );
  OAI222 U3811 ( .A(n628), .B(n10966), .C(n604), .D(n11235), .Q(n10236) );
  OAI222 U3812 ( .A(n580), .B(n10964), .C(n556), .D(n11234), .Q(n10235) );
  OAI222 U3816 ( .A(n5524), .B(n10962), .C(n5500), .D(n11233), .Q(n10250) );
  OAI222 U3817 ( .A(n5476), .B(n10960), .C(n5452), .D(n11232), .Q(n10249) );
  OAI222 U3818 ( .A(n5428), .B(n10958), .C(n5404), .D(n11231), .Q(n10248) );
  OAI222 U3819 ( .A(n5380), .B(n10956), .C(n5356), .D(n11230), .Q(n10247) );
  OAI222 U3821 ( .A(n5716), .B(n10954), .C(n5692), .D(n11229), .Q(n10254) );
  OAI222 U3822 ( .A(n5668), .B(n10952), .C(n5644), .D(n11228), .Q(n10253) );
  OAI222 U3823 ( .A(n5620), .B(n10950), .C(n5596), .D(n11227), .Q(n10252) );
  OAI222 U3824 ( .A(n5572), .B(n10948), .C(n5548), .D(n11226), .Q(n10251) );
  OAI222 U3826 ( .A(n5908), .B(n10946), .C(n5884), .D(n11225), .Q(n10258) );
  OAI222 U3827 ( .A(n5860), .B(n10944), .C(n5836), .D(n11224), .Q(n10257) );
  OAI222 U3828 ( .A(n5812), .B(n10942), .C(n5788), .D(n11223), .Q(n10256) );
  OAI222 U3829 ( .A(n5764), .B(n10940), .C(n5740), .D(n11222), .Q(n10255) );
  OAI222 U3831 ( .A(n6100), .B(n10938), .C(n6076), .D(n11221), .Q(n10262) );
  OAI222 U3832 ( .A(n6052), .B(n10936), .C(n6028), .D(n11220), .Q(n10261) );
  OAI222 U3833 ( .A(n6004), .B(n10934), .C(n5980), .D(n11219), .Q(n10260) );
  OAI222 U3834 ( .A(n5956), .B(n10932), .C(n5932), .D(n11218), .Q(n10259) );
  OAI222 U3837 ( .A(n4756), .B(n10930), .C(n4732), .D(n11217), .Q(n10270) );
  OAI222 U3838 ( .A(n4708), .B(n10928), .C(n4684), .D(n11216), .Q(n10269) );
  OAI222 U3839 ( .A(n4660), .B(n10926), .C(n4636), .D(n11215), .Q(n10268) );
  OAI222 U3840 ( .A(n4612), .B(n10924), .C(n4588), .D(n11214), .Q(n10267) );
  OAI222 U3842 ( .A(n4948), .B(n10922), .C(n4924), .D(n11213), .Q(n10274) );
  OAI222 U3843 ( .A(n4900), .B(n10920), .C(n4876), .D(n11212), .Q(n10273) );
  OAI222 U3844 ( .A(n4852), .B(n10918), .C(n4828), .D(n11211), .Q(n10272) );
  OAI222 U3845 ( .A(n4804), .B(n10916), .C(n4780), .D(n11210), .Q(n10271) );
  OAI222 U3847 ( .A(n5140), .B(n10914), .C(n5116), .D(n11209), .Q(n10278) );
  OAI222 U3848 ( .A(n5092), .B(n10912), .C(n5068), .D(n11208), .Q(n10277) );
  OAI222 U3849 ( .A(n5044), .B(n10910), .C(n5020), .D(n11207), .Q(n10276) );
  OAI222 U3850 ( .A(n4996), .B(n10908), .C(n4972), .D(n11206), .Q(n10275) );
  OAI222 U3852 ( .A(n5332), .B(n10906), .C(n5308), .D(n11205), .Q(n10282) );
  OAI222 U3853 ( .A(n5284), .B(n10904), .C(n5260), .D(n11204), .Q(n10281) );
  OAI222 U3854 ( .A(n5236), .B(n10902), .C(n5212), .D(n11203), .Q(n10280) );
  OAI222 U3855 ( .A(n5188), .B(n10900), .C(n5164), .D(n11202), .Q(n10279) );
  OAI222 U3858 ( .A(n3988), .B(n10898), .C(n3964), .D(n11201), .Q(n10290) );
  OAI222 U3859 ( .A(n3940), .B(n10896), .C(n3916), .D(n11200), .Q(n10289) );
  OAI222 U3860 ( .A(n3892), .B(n10894), .C(n3868), .D(n11199), .Q(n10288) );
  OAI222 U3861 ( .A(n3844), .B(n10892), .C(n3820), .D(n11198), .Q(n10287) );
  OAI222 U3863 ( .A(n4180), .B(n10890), .C(n4156), .D(n11197), .Q(n10294) );
  OAI222 U3864 ( .A(n4132), .B(n10888), .C(n4108), .D(n11196), .Q(n10293) );
  OAI222 U3865 ( .A(n4084), .B(n10886), .C(n4060), .D(n11195), .Q(n10292) );
  OAI222 U3866 ( .A(n4036), .B(n10884), .C(n4012), .D(n11194), .Q(n10291) );
  OAI222 U3868 ( .A(n4372), .B(n10882), .C(n4348), .D(n11193), .Q(n10298) );
  OAI222 U3869 ( .A(n4324), .B(n6192), .C(n4300), .D(n11192), .Q(n10297) );
  OAI222 U3870 ( .A(n4276), .B(n6190), .C(n4252), .D(n11191), .Q(n10296) );
  OAI222 U3871 ( .A(n4228), .B(n6188), .C(n4204), .D(n11190), .Q(n10295) );
  OAI222 U3873 ( .A(n4564), .B(n6186), .C(n4540), .D(n11189), .Q(n10302) );
  OAI222 U3874 ( .A(n4516), .B(n6184), .C(n4492), .D(n11188), .Q(n10301) );
  OAI222 U3875 ( .A(n4468), .B(n6182), .C(n4444), .D(n11187), .Q(n10300) );
  OAI222 U3876 ( .A(n4420), .B(n6180), .C(n4396), .D(n11186), .Q(n10299) );
  OAI222 U3879 ( .A(n3220), .B(n6178), .C(n3196), .D(n11185), .Q(n10310) );
  OAI222 U3880 ( .A(n3172), .B(n6176), .C(n3148), .D(n11184), .Q(n10309) );
  OAI222 U3881 ( .A(n3124), .B(n6174), .C(n3100), .D(n11183), .Q(n10308) );
  OAI222 U3882 ( .A(n3076), .B(n6172), .C(n3052), .D(n11182), .Q(n10307) );
  OAI222 U3884 ( .A(n3412), .B(n6170), .C(n3388), .D(n11181), .Q(n10314) );
  OAI222 U3885 ( .A(n3364), .B(n6168), .C(n3340), .D(n11180), .Q(n10313) );
  OAI222 U3886 ( .A(n3316), .B(n6166), .C(n3292), .D(n11179), .Q(n10312) );
  OAI222 U3887 ( .A(n3268), .B(n6164), .C(n3244), .D(n11178), .Q(n10311) );
  OAI222 U3889 ( .A(n3604), .B(n6162), .C(n3580), .D(n11177), .Q(n10318) );
  OAI222 U3890 ( .A(n3556), .B(n6160), .C(n3532), .D(n11176), .Q(n10317) );
  OAI222 U3891 ( .A(n3508), .B(n6158), .C(n3484), .D(n11175), .Q(n10316) );
  OAI222 U3892 ( .A(n3460), .B(n6156), .C(n3436), .D(n11174), .Q(n10315) );
  OAI222 U3894 ( .A(n3796), .B(n6154), .C(n3772), .D(n11173), .Q(n10322) );
  OAI222 U3895 ( .A(n3748), .B(n6152), .C(n3724), .D(n11172), .Q(n10321) );
  OAI222 U3896 ( .A(n3700), .B(n6150), .C(n3676), .D(n11171), .Q(n10320) );
  OAI222 U3897 ( .A(n3652), .B(n6148), .C(n3628), .D(n11170), .Q(n10319) );
  OAI222 U3902 ( .A(n2451), .B(n11090), .C(n2427), .D(n11297), .Q(n10336) );
  OAI222 U3903 ( .A(n2403), .B(n11088), .C(n2379), .D(n11296), .Q(n10335) );
  OAI222 U3904 ( .A(n2355), .B(n11086), .C(n2331), .D(n11295), .Q(n10334) );
  OAI222 U3905 ( .A(n2307), .B(n11084), .C(n2283), .D(n11294), .Q(n10333) );
  OAI222 U3907 ( .A(n2643), .B(n11082), .C(n2619), .D(n11293), .Q(n10340) );
  OAI222 U3908 ( .A(n2595), .B(n11080), .C(n2571), .D(n11292), .Q(n10339) );
  OAI222 U3909 ( .A(n2547), .B(n11078), .C(n2523), .D(n11291), .Q(n10338) );
  OAI222 U3910 ( .A(n2499), .B(n11076), .C(n2475), .D(n11290), .Q(n10337) );
  OAI222 U3912 ( .A(n2835), .B(n11074), .C(n2811), .D(n11289), .Q(n10344) );
  OAI222 U3913 ( .A(n2787), .B(n11072), .C(n2763), .D(n11288), .Q(n10343) );
  OAI222 U3914 ( .A(n2739), .B(n11070), .C(n2715), .D(n11287), .Q(n10342) );
  OAI222 U3915 ( .A(n2691), .B(n11068), .C(n2667), .D(n11286), .Q(n10341) );
  OAI222 U3917 ( .A(n3027), .B(n11066), .C(n3003), .D(n11285), .Q(n10348) );
  OAI222 U3918 ( .A(n2979), .B(n11064), .C(n2955), .D(n11284), .Q(n10347) );
  OAI222 U3919 ( .A(n2931), .B(n11062), .C(n2907), .D(n11283), .Q(n10346) );
  OAI222 U3920 ( .A(n2883), .B(n11060), .C(n2859), .D(n11282), .Q(n10345) );
  OAI222 U3923 ( .A(n1683), .B(n11058), .C(n1659), .D(n11281), .Q(n10356) );
  OAI222 U3924 ( .A(n1635), .B(n11056), .C(n1611), .D(n11280), .Q(n10355) );
  OAI222 U3925 ( .A(n1587), .B(n11054), .C(n1563), .D(n11279), .Q(n10354) );
  OAI222 U3926 ( .A(n1539), .B(n11052), .C(n1515), .D(n11278), .Q(n10353) );
  OAI222 U3928 ( .A(n1875), .B(n11050), .C(n1851), .D(n11277), .Q(n10360) );
  OAI222 U3929 ( .A(n1827), .B(n11048), .C(n1803), .D(n11276), .Q(n10359) );
  OAI222 U3930 ( .A(n1779), .B(n11046), .C(n1755), .D(n11275), .Q(n10358) );
  OAI222 U3931 ( .A(n1731), .B(n11044), .C(n1707), .D(n11274), .Q(n10357) );
  OAI222 U3933 ( .A(n2067), .B(n11042), .C(n2043), .D(n11273), .Q(n10364) );
  OAI222 U3934 ( .A(n2019), .B(n11040), .C(n1995), .D(n11272), .Q(n10363) );
  OAI222 U3935 ( .A(n1971), .B(n11038), .C(n1947), .D(n11271), .Q(n10362) );
  OAI222 U3936 ( .A(n1923), .B(n11036), .C(n1899), .D(n11270), .Q(n10361) );
  OAI222 U3938 ( .A(n2259), .B(n11034), .C(n2235), .D(n11269), .Q(n10368) );
  OAI222 U3939 ( .A(n2211), .B(n11032), .C(n2187), .D(n11268), .Q(n10367) );
  OAI222 U3940 ( .A(n2163), .B(n11030), .C(n2139), .D(n11267), .Q(n10366) );
  OAI222 U3941 ( .A(n2115), .B(n11028), .C(n2091), .D(n11266), .Q(n10365) );
  OAI222 U3944 ( .A(n915), .B(n11026), .C(n891), .D(n11265), .Q(n10376) );
  OAI222 U3945 ( .A(n867), .B(n11024), .C(n843), .D(n11264), .Q(n10375) );
  OAI222 U3946 ( .A(n819), .B(n11022), .C(n795), .D(n11263), .Q(n10374) );
  OAI222 U3947 ( .A(n771), .B(n11020), .C(n747), .D(n11262), .Q(n10373) );
  OAI222 U3949 ( .A(n1107), .B(n11018), .C(n1083), .D(n11261), .Q(n10380) );
  OAI222 U3950 ( .A(n1059), .B(n11016), .C(n1035), .D(n11260), .Q(n10379) );
  OAI222 U3951 ( .A(n1011), .B(n11014), .C(n987), .D(n11259), .Q(n10378) );
  OAI222 U3952 ( .A(n963), .B(n11012), .C(n939), .D(n11258), .Q(n10377) );
  OAI222 U3954 ( .A(n1299), .B(n11010), .C(n1275), .D(n11257), .Q(n10384) );
  OAI222 U3955 ( .A(n1251), .B(n11008), .C(n1227), .D(n11256), .Q(n10383) );
  OAI222 U3956 ( .A(n1203), .B(n11006), .C(n1179), .D(n11255), .Q(n10382) );
  OAI222 U3957 ( .A(n1155), .B(n11004), .C(n1131), .D(n11254), .Q(n10381) );
  OAI222 U3959 ( .A(n1491), .B(n11002), .C(n1467), .D(n11253), .Q(n10388) );
  OAI222 U3960 ( .A(n1443), .B(n11000), .C(n1419), .D(n11252), .Q(n10387) );
  OAI222 U3961 ( .A(n1395), .B(n10998), .C(n1371), .D(n11251), .Q(n10386) );
  OAI222 U3962 ( .A(n1347), .B(n10996), .C(n1323), .D(n11250), .Q(n10385) );
  OAI222 U3965 ( .A(n147), .B(n10994), .C(n123), .D(n11249), .Q(n10396) );
  OAI222 U3966 ( .A(n99), .B(n10992), .C(n75), .D(n11248), .Q(n10395) );
  OAI222 U3967 ( .A(n51), .B(n10990), .C(n27), .D(n11247), .Q(n10394) );
  OAI222 U3968 ( .A(n3), .B(n10988), .C(n6123), .D(n11246), .Q(n10393) );
  OAI222 U3970 ( .A(n339), .B(n10986), .C(n315), .D(n11245), .Q(n10400) );
  OAI222 U3971 ( .A(n291), .B(n10984), .C(n267), .D(n11244), .Q(n10399) );
  OAI222 U3972 ( .A(n243), .B(n10982), .C(n219), .D(n11243), .Q(n10398) );
  OAI222 U3973 ( .A(n195), .B(n10980), .C(n171), .D(n11242), .Q(n10397) );
  OAI222 U3975 ( .A(n531), .B(n10978), .C(n507), .D(n11241), .Q(n10404) );
  OAI222 U3976 ( .A(n483), .B(n10976), .C(n459), .D(n11240), .Q(n10403) );
  OAI222 U3977 ( .A(n435), .B(n10974), .C(n411), .D(n11239), .Q(n10402) );
  OAI222 U3978 ( .A(n387), .B(n10972), .C(n363), .D(n11238), .Q(n10401) );
  OAI222 U3980 ( .A(n723), .B(n10970), .C(n699), .D(n11237), .Q(n10408) );
  OAI222 U3981 ( .A(n675), .B(n10968), .C(n651), .D(n11236), .Q(n10407) );
  OAI222 U3982 ( .A(n627), .B(n10966), .C(n603), .D(n11235), .Q(n10406) );
  OAI222 U3983 ( .A(n579), .B(n10964), .C(n555), .D(n11234), .Q(n10405) );
  OAI222 U3987 ( .A(n5523), .B(n10962), .C(n5499), .D(n11233), .Q(n10420) );
  OAI222 U3988 ( .A(n5475), .B(n10960), .C(n5451), .D(n11232), .Q(n10419) );
  OAI222 U3989 ( .A(n5427), .B(n10958), .C(n5403), .D(n11231), .Q(n10418) );
  OAI222 U3990 ( .A(n5379), .B(n10956), .C(n5355), .D(n11230), .Q(n10417) );
  OAI222 U3992 ( .A(n5715), .B(n10954), .C(n5691), .D(n11229), .Q(n10424) );
  OAI222 U3993 ( .A(n5667), .B(n10952), .C(n5643), .D(n11228), .Q(n10423) );
  OAI222 U3994 ( .A(n5619), .B(n10950), .C(n5595), .D(n11227), .Q(n10422) );
  OAI222 U3995 ( .A(n5571), .B(n10948), .C(n5547), .D(n11226), .Q(n10421) );
  OAI222 U3997 ( .A(n5907), .B(n10946), .C(n5883), .D(n11225), .Q(n10428) );
  OAI222 U3998 ( .A(n5859), .B(n10944), .C(n5835), .D(n11224), .Q(n10427) );
  OAI222 U3999 ( .A(n5811), .B(n10942), .C(n5787), .D(n11223), .Q(n10426) );
  OAI222 U4000 ( .A(n5763), .B(n10940), .C(n5739), .D(n11222), .Q(n10425) );
  OAI222 U4002 ( .A(n6099), .B(n10938), .C(n6075), .D(n11221), .Q(n10432) );
  OAI222 U4003 ( .A(n6051), .B(n10936), .C(n6027), .D(n11220), .Q(n10431) );
  OAI222 U4004 ( .A(n6003), .B(n10934), .C(n5979), .D(n11219), .Q(n10430) );
  OAI222 U4005 ( .A(n5955), .B(n10932), .C(n5931), .D(n11218), .Q(n10429) );
  OAI222 U4008 ( .A(n4755), .B(n10930), .C(n4731), .D(n11217), .Q(n10440) );
  OAI222 U4009 ( .A(n4707), .B(n10928), .C(n4683), .D(n11216), .Q(n10439) );
  OAI222 U4010 ( .A(n4659), .B(n10926), .C(n4635), .D(n11215), .Q(n10438) );
  OAI222 U4011 ( .A(n4611), .B(n10924), .C(n4587), .D(n11214), .Q(n10437) );
  OAI222 U4013 ( .A(n4947), .B(n10922), .C(n4923), .D(n11213), .Q(n10444) );
  OAI222 U4014 ( .A(n4899), .B(n10920), .C(n4875), .D(n11212), .Q(n10443) );
  OAI222 U4015 ( .A(n4851), .B(n10918), .C(n4827), .D(n11211), .Q(n10442) );
  OAI222 U4016 ( .A(n4803), .B(n10916), .C(n4779), .D(n11210), .Q(n10441) );
  OAI222 U4018 ( .A(n5139), .B(n10914), .C(n5115), .D(n11209), .Q(n10448) );
  OAI222 U4019 ( .A(n5091), .B(n10912), .C(n5067), .D(n11208), .Q(n10447) );
  OAI222 U4020 ( .A(n5043), .B(n10910), .C(n5019), .D(n11207), .Q(n10446) );
  OAI222 U4021 ( .A(n4995), .B(n10908), .C(n4971), .D(n11206), .Q(n10445) );
  OAI222 U4023 ( .A(n5331), .B(n10906), .C(n5307), .D(n11205), .Q(n10452) );
  OAI222 U4024 ( .A(n5283), .B(n10904), .C(n5259), .D(n11204), .Q(n10451) );
  OAI222 U4025 ( .A(n5235), .B(n10902), .C(n5211), .D(n11203), .Q(n10450) );
  OAI222 U4026 ( .A(n5187), .B(n10900), .C(n5163), .D(n11202), .Q(n10449) );
  OAI222 U4029 ( .A(n3987), .B(n10898), .C(n3963), .D(n11201), .Q(n10460) );
  OAI222 U4030 ( .A(n3939), .B(n10896), .C(n3915), .D(n11200), .Q(n10459) );
  OAI222 U4031 ( .A(n3891), .B(n10894), .C(n3867), .D(n11199), .Q(n10458) );
  OAI222 U4032 ( .A(n3843), .B(n10892), .C(n3819), .D(n11198), .Q(n10457) );
  OAI222 U4034 ( .A(n4179), .B(n10890), .C(n4155), .D(n11197), .Q(n10464) );
  OAI222 U4035 ( .A(n4131), .B(n10888), .C(n4107), .D(n11196), .Q(n10463) );
  OAI222 U4036 ( .A(n4083), .B(n10886), .C(n4059), .D(n11195), .Q(n10462) );
  OAI222 U4037 ( .A(n4035), .B(n10884), .C(n4011), .D(n11194), .Q(n10461) );
  OAI222 U4039 ( .A(n4371), .B(n10882), .C(n4347), .D(n11193), .Q(n10468) );
  OAI222 U4040 ( .A(n4323), .B(n6192), .C(n4299), .D(n11192), .Q(n10467) );
  OAI222 U4041 ( .A(n4275), .B(n6190), .C(n4251), .D(n11191), .Q(n10466) );
  OAI222 U4042 ( .A(n4227), .B(n6188), .C(n4203), .D(n11190), .Q(n10465) );
  OAI222 U4044 ( .A(n4563), .B(n6186), .C(n4539), .D(n11189), .Q(n10472) );
  OAI222 U4045 ( .A(n4515), .B(n6184), .C(n4491), .D(n11188), .Q(n10471) );
  OAI222 U4046 ( .A(n4467), .B(n6182), .C(n4443), .D(n11187), .Q(n10470) );
  OAI222 U4047 ( .A(n4419), .B(n6180), .C(n4395), .D(n11186), .Q(n10469) );
  OAI222 U4050 ( .A(n3219), .B(n6178), .C(n3195), .D(n11185), .Q(n10480) );
  OAI222 U4051 ( .A(n3171), .B(n6176), .C(n3147), .D(n11184), .Q(n10479) );
  OAI222 U4052 ( .A(n3123), .B(n6174), .C(n3099), .D(n11183), .Q(n10478) );
  OAI222 U4053 ( .A(n3075), .B(n6172), .C(n3051), .D(n11182), .Q(n10477) );
  OAI222 U4055 ( .A(n3411), .B(n6170), .C(n3387), .D(n11181), .Q(n10484) );
  OAI222 U4056 ( .A(n3363), .B(n6168), .C(n3339), .D(n11180), .Q(n10483) );
  OAI222 U4057 ( .A(n3315), .B(n6166), .C(n3291), .D(n11179), .Q(n10482) );
  OAI222 U4058 ( .A(n3267), .B(n6164), .C(n3243), .D(n11178), .Q(n10481) );
  OAI222 U4060 ( .A(n3603), .B(n6162), .C(n3579), .D(n11177), .Q(n10488) );
  OAI222 U4061 ( .A(n3555), .B(n6160), .C(n3531), .D(n11176), .Q(n10487) );
  OAI222 U4062 ( .A(n3507), .B(n6158), .C(n3483), .D(n11175), .Q(n10486) );
  OAI222 U4063 ( .A(n3459), .B(n6156), .C(n3435), .D(n11174), .Q(n10485) );
  OAI222 U4065 ( .A(n3795), .B(n6154), .C(n3771), .D(n11173), .Q(n10492) );
  OAI222 U4066 ( .A(n3747), .B(n6152), .C(n3723), .D(n11172), .Q(n10491) );
  OAI222 U4067 ( .A(n3699), .B(n6150), .C(n3675), .D(n11171), .Q(n10490) );
  OAI222 U4068 ( .A(n3651), .B(n6148), .C(n3627), .D(n11170), .Q(n10489) );
  OAI222 U4073 ( .A(n2450), .B(n11090), .C(n2426), .D(n11297), .Q(n10506) );
  OAI222 U4074 ( .A(n2402), .B(n11088), .C(n2378), .D(n11296), .Q(n10505) );
  OAI222 U4075 ( .A(n2354), .B(n11086), .C(n2330), .D(n11295), .Q(n10504) );
  OAI222 U4076 ( .A(n2306), .B(n11084), .C(n2282), .D(n11294), .Q(n10503) );
  OAI222 U4078 ( .A(n2642), .B(n11082), .C(n2618), .D(n11293), .Q(n10510) );
  OAI222 U4079 ( .A(n2594), .B(n11080), .C(n2570), .D(n11292), .Q(n10509) );
  OAI222 U4080 ( .A(n2546), .B(n11078), .C(n2522), .D(n11291), .Q(n10508) );
  OAI222 U4081 ( .A(n2498), .B(n11076), .C(n2474), .D(n11290), .Q(n10507) );
  OAI222 U4083 ( .A(n2834), .B(n11074), .C(n2810), .D(n11289), .Q(n10514) );
  OAI222 U4084 ( .A(n2786), .B(n11072), .C(n2762), .D(n11288), .Q(n10513) );
  OAI222 U4085 ( .A(n2738), .B(n11070), .C(n2714), .D(n11287), .Q(n10512) );
  OAI222 U4086 ( .A(n2690), .B(n11068), .C(n2666), .D(n11286), .Q(n10511) );
  OAI222 U4088 ( .A(n3026), .B(n11066), .C(n3002), .D(n11285), .Q(n10518) );
  OAI222 U4089 ( .A(n2978), .B(n11064), .C(n2954), .D(n11284), .Q(n10517) );
  OAI222 U4090 ( .A(n2930), .B(n11062), .C(n2906), .D(n11283), .Q(n10516) );
  OAI222 U4091 ( .A(n2882), .B(n11060), .C(n2858), .D(n11282), .Q(n10515) );
  OAI222 U4094 ( .A(n1682), .B(n11058), .C(n1658), .D(n11281), .Q(n10526) );
  OAI222 U4095 ( .A(n1634), .B(n11056), .C(n1610), .D(n11280), .Q(n10525) );
  OAI222 U4096 ( .A(n1586), .B(n11054), .C(n1562), .D(n11279), .Q(n10524) );
  OAI222 U4097 ( .A(n1538), .B(n11052), .C(n1514), .D(n11278), .Q(n10523) );
  OAI222 U4099 ( .A(n1874), .B(n11050), .C(n1850), .D(n11277), .Q(n10530) );
  OAI222 U4100 ( .A(n1826), .B(n11048), .C(n1802), .D(n11276), .Q(n10529) );
  OAI222 U4101 ( .A(n1778), .B(n11046), .C(n1754), .D(n11275), .Q(n10528) );
  OAI222 U4102 ( .A(n1730), .B(n11044), .C(n1706), .D(n11274), .Q(n10527) );
  OAI222 U4104 ( .A(n2066), .B(n11042), .C(n2042), .D(n11273), .Q(n10534) );
  OAI222 U4105 ( .A(n2018), .B(n11040), .C(n1994), .D(n11272), .Q(n10533) );
  OAI222 U4106 ( .A(n1970), .B(n11038), .C(n1946), .D(n11271), .Q(n10532) );
  OAI222 U4107 ( .A(n1922), .B(n11036), .C(n1898), .D(n11270), .Q(n10531) );
  OAI222 U4109 ( .A(n2258), .B(n11034), .C(n2234), .D(n11269), .Q(n10538) );
  OAI222 U4110 ( .A(n2210), .B(n11032), .C(n2186), .D(n11268), .Q(n10537) );
  OAI222 U4111 ( .A(n2162), .B(n11030), .C(n2138), .D(n11267), .Q(n10536) );
  OAI222 U4112 ( .A(n2114), .B(n11028), .C(n2090), .D(n11266), .Q(n10535) );
  OAI222 U4115 ( .A(n914), .B(n11026), .C(n890), .D(n11265), .Q(n10546) );
  OAI222 U4116 ( .A(n866), .B(n11024), .C(n842), .D(n11264), .Q(n10545) );
  OAI222 U4117 ( .A(n818), .B(n11022), .C(n794), .D(n11263), .Q(n10544) );
  OAI222 U4118 ( .A(n770), .B(n11020), .C(n746), .D(n11262), .Q(n10543) );
  OAI222 U4120 ( .A(n1106), .B(n11018), .C(n1082), .D(n11261), .Q(n10550) );
  OAI222 U4121 ( .A(n1058), .B(n11016), .C(n1034), .D(n11260), .Q(n10549) );
  OAI222 U4122 ( .A(n1010), .B(n11014), .C(n986), .D(n11259), .Q(n10548) );
  OAI222 U4123 ( .A(n962), .B(n11012), .C(n938), .D(n11258), .Q(n10547) );
  OAI222 U4125 ( .A(n1298), .B(n11010), .C(n1274), .D(n11257), .Q(n10554) );
  OAI222 U4126 ( .A(n1250), .B(n11008), .C(n1226), .D(n11256), .Q(n10553) );
  OAI222 U4127 ( .A(n1202), .B(n11006), .C(n1178), .D(n11255), .Q(n10552) );
  OAI222 U4128 ( .A(n1154), .B(n11004), .C(n1130), .D(n11254), .Q(n10551) );
  OAI222 U4130 ( .A(n1490), .B(n11002), .C(n1466), .D(n11253), .Q(n10558) );
  OAI222 U4131 ( .A(n1442), .B(n11000), .C(n1418), .D(n11252), .Q(n10557) );
  OAI222 U4132 ( .A(n1394), .B(n10998), .C(n1370), .D(n11251), .Q(n10556) );
  OAI222 U4133 ( .A(n1346), .B(n10996), .C(n1322), .D(n11250), .Q(n10555) );
  OAI222 U4136 ( .A(n146), .B(n10994), .C(n122), .D(n11249), .Q(n10566) );
  OAI222 U4137 ( .A(n98), .B(n10992), .C(n74), .D(n11248), .Q(n10565) );
  OAI222 U4138 ( .A(n50), .B(n10990), .C(n26), .D(n11247), .Q(n10564) );
  OAI222 U4139 ( .A(n2), .B(n10988), .C(n6122), .D(n11246), .Q(n10563) );
  OAI222 U4141 ( .A(n338), .B(n10986), .C(n314), .D(n11245), .Q(n10570) );
  OAI222 U4142 ( .A(n290), .B(n10984), .C(n266), .D(n11244), .Q(n10569) );
  OAI222 U4143 ( .A(n242), .B(n10982), .C(n218), .D(n11243), .Q(n10568) );
  OAI222 U4144 ( .A(n194), .B(n10980), .C(n170), .D(n11242), .Q(n10567) );
  OAI222 U4146 ( .A(n530), .B(n10978), .C(n506), .D(n11241), .Q(n10574) );
  OAI222 U4147 ( .A(n482), .B(n10976), .C(n458), .D(n11240), .Q(n10573) );
  OAI222 U4148 ( .A(n434), .B(n10974), .C(n410), .D(n11239), .Q(n10572) );
  OAI222 U4149 ( .A(n386), .B(n10972), .C(n362), .D(n11238), .Q(n10571) );
  OAI222 U4151 ( .A(n722), .B(n10970), .C(n698), .D(n11237), .Q(n10578) );
  OAI222 U4152 ( .A(n674), .B(n10968), .C(n650), .D(n11236), .Q(n10577) );
  OAI222 U4153 ( .A(n626), .B(n10966), .C(n602), .D(n11235), .Q(n10576) );
  OAI222 U4154 ( .A(n578), .B(n10964), .C(n554), .D(n11234), .Q(n10575) );
  OAI222 U4158 ( .A(n5522), .B(n10962), .C(n5498), .D(n11233), .Q(n10590) );
  OAI222 U4159 ( .A(n5474), .B(n10960), .C(n5450), .D(n11232), .Q(n10589) );
  OAI222 U4160 ( .A(n5426), .B(n10958), .C(n5402), .D(n11231), .Q(n10588) );
  OAI222 U4161 ( .A(n5378), .B(n10956), .C(n5354), .D(n11230), .Q(n10587) );
  OAI222 U4163 ( .A(n5714), .B(n10954), .C(n5690), .D(n11229), .Q(n10594) );
  OAI222 U4164 ( .A(n5666), .B(n10952), .C(n5642), .D(n11228), .Q(n10593) );
  OAI222 U4165 ( .A(n5618), .B(n10950), .C(n5594), .D(n11227), .Q(n10592) );
  OAI222 U4166 ( .A(n5570), .B(n10948), .C(n5546), .D(n11226), .Q(n10591) );
  OAI222 U4168 ( .A(n5906), .B(n10946), .C(n5882), .D(n11225), .Q(n10598) );
  OAI222 U4169 ( .A(n5858), .B(n10944), .C(n5834), .D(n11224), .Q(n10597) );
  OAI222 U4170 ( .A(n5810), .B(n10942), .C(n5786), .D(n11223), .Q(n10596) );
  OAI222 U4171 ( .A(n5762), .B(n10940), .C(n5738), .D(n11222), .Q(n10595) );
  OAI222 U4173 ( .A(n6098), .B(n10938), .C(n6074), .D(n11221), .Q(n10602) );
  OAI222 U4174 ( .A(n6050), .B(n10936), .C(n6026), .D(n11220), .Q(n10601) );
  OAI222 U4175 ( .A(n6002), .B(n10934), .C(n5978), .D(n11219), .Q(n10600) );
  OAI222 U4176 ( .A(n5954), .B(n10932), .C(n5930), .D(n11218), .Q(n10599) );
  OAI222 U4179 ( .A(n4754), .B(n10930), .C(n4730), .D(n11217), .Q(n10610) );
  OAI222 U4180 ( .A(n4706), .B(n10928), .C(n4682), .D(n11216), .Q(n10609) );
  OAI222 U4181 ( .A(n4658), .B(n10926), .C(n4634), .D(n11215), .Q(n10608) );
  OAI222 U4182 ( .A(n4610), .B(n10924), .C(n4586), .D(n11214), .Q(n10607) );
  OAI222 U4184 ( .A(n4946), .B(n10922), .C(n4922), .D(n11213), .Q(n10614) );
  OAI222 U4185 ( .A(n4898), .B(n10920), .C(n4874), .D(n11212), .Q(n10613) );
  OAI222 U4186 ( .A(n4850), .B(n10918), .C(n4826), .D(n11211), .Q(n10612) );
  OAI222 U4187 ( .A(n4802), .B(n10916), .C(n4778), .D(n11210), .Q(n10611) );
  OAI222 U4189 ( .A(n5138), .B(n10914), .C(n5114), .D(n11209), .Q(n10618) );
  OAI222 U4190 ( .A(n5090), .B(n10912), .C(n5066), .D(n11208), .Q(n10617) );
  OAI222 U4191 ( .A(n5042), .B(n10910), .C(n5018), .D(n11207), .Q(n10616) );
  OAI222 U4192 ( .A(n4994), .B(n10908), .C(n4970), .D(n11206), .Q(n10615) );
  OAI222 U4194 ( .A(n5330), .B(n10906), .C(n5306), .D(n11205), .Q(n10622) );
  OAI222 U4195 ( .A(n5282), .B(n10904), .C(n5258), .D(n11204), .Q(n10621) );
  OAI222 U4196 ( .A(n5234), .B(n10902), .C(n5210), .D(n11203), .Q(n10620) );
  OAI222 U4197 ( .A(n5186), .B(n10900), .C(n5162), .D(n11202), .Q(n10619) );
  OAI222 U4200 ( .A(n3986), .B(n10898), .C(n3962), .D(n11201), .Q(n10630) );
  OAI222 U4201 ( .A(n3938), .B(n10896), .C(n3914), .D(n11200), .Q(n10629) );
  OAI222 U4202 ( .A(n3890), .B(n10894), .C(n3866), .D(n11199), .Q(n10628) );
  OAI222 U4203 ( .A(n3842), .B(n10892), .C(n3818), .D(n11198), .Q(n10627) );
  OAI222 U4205 ( .A(n4178), .B(n10890), .C(n4154), .D(n11197), .Q(n10634) );
  OAI222 U4206 ( .A(n4130), .B(n10888), .C(n4106), .D(n11196), .Q(n10633) );
  OAI222 U4207 ( .A(n4082), .B(n10886), .C(n4058), .D(n11195), .Q(n10632) );
  OAI222 U4208 ( .A(n4034), .B(n10884), .C(n4010), .D(n11194), .Q(n10631) );
  OAI222 U4210 ( .A(n4370), .B(n10882), .C(n4346), .D(n11193), .Q(n10638) );
  OAI222 U4211 ( .A(n4322), .B(n6192), .C(n4298), .D(n11192), .Q(n10637) );
  OAI222 U4212 ( .A(n4274), .B(n6190), .C(n4250), .D(n11191), .Q(n10636) );
  OAI222 U4213 ( .A(n4226), .B(n6188), .C(n4202), .D(n11190), .Q(n10635) );
  OAI222 U4215 ( .A(n4562), .B(n6186), .C(n4538), .D(n11189), .Q(n10642) );
  OAI222 U4216 ( .A(n4514), .B(n6184), .C(n4490), .D(n11188), .Q(n10641) );
  OAI222 U4217 ( .A(n4466), .B(n6182), .C(n4442), .D(n11187), .Q(n10640) );
  OAI222 U4218 ( .A(n4418), .B(n6180), .C(n4394), .D(n11186), .Q(n10639) );
  OAI222 U4221 ( .A(n3218), .B(n6178), .C(n3194), .D(n11185), .Q(n10650) );
  OAI222 U4222 ( .A(n3170), .B(n6176), .C(n3146), .D(n11184), .Q(n10649) );
  OAI222 U4223 ( .A(n3122), .B(n6174), .C(n3098), .D(n11183), .Q(n10648) );
  OAI222 U4224 ( .A(n3074), .B(n6172), .C(n3050), .D(n11182), .Q(n10647) );
  OAI222 U4226 ( .A(n3410), .B(n6170), .C(n3386), .D(n11181), .Q(n10654) );
  OAI222 U4227 ( .A(n3362), .B(n6168), .C(n3338), .D(n11180), .Q(n10653) );
  OAI222 U4228 ( .A(n3314), .B(n6166), .C(n3290), .D(n11179), .Q(n10652) );
  OAI222 U4229 ( .A(n3266), .B(n6164), .C(n3242), .D(n11178), .Q(n10651) );
  OAI222 U4231 ( .A(n3602), .B(n6162), .C(n3578), .D(n11177), .Q(n10658) );
  OAI222 U4232 ( .A(n3554), .B(n6160), .C(n3530), .D(n11176), .Q(n10657) );
  OAI222 U4233 ( .A(n3506), .B(n6158), .C(n3482), .D(n11175), .Q(n10656) );
  OAI222 U4234 ( .A(n3458), .B(n6156), .C(n3434), .D(n11174), .Q(n10655) );
  OAI222 U4236 ( .A(n3794), .B(n6154), .C(n3770), .D(n11173), .Q(n10662) );
  OAI222 U4237 ( .A(n3746), .B(n6152), .C(n3722), .D(n11172), .Q(n10661) );
  OAI222 U4238 ( .A(n3698), .B(n6150), .C(n3674), .D(n11171), .Q(n10660) );
  OAI222 U4239 ( .A(n3650), .B(n6148), .C(n3626), .D(n11170), .Q(n10659) );
  OAI222 U4244 ( .A(n2449), .B(n11090), .C(n2425), .D(n11297), .Q(n10676) );
  OAI222 U4247 ( .A(n2401), .B(n11088), .C(n2377), .D(n11296), .Q(n10675) );
  OAI222 U4250 ( .A(n2353), .B(n11086), .C(n2329), .D(n11295), .Q(n10674) );
  OAI222 U4253 ( .A(n2305), .B(n11084), .C(n2281), .D(n11294), .Q(n10673) );
  OAI222 U4257 ( .A(n2641), .B(n11082), .C(n2617), .D(n11293), .Q(n10680) );
  OAI222 U4260 ( .A(n2593), .B(n11080), .C(n2569), .D(n11292), .Q(n10679) );
  OAI222 U4263 ( .A(n2545), .B(n11078), .C(n2521), .D(n11291), .Q(n10678) );
  OAI222 U4266 ( .A(n2497), .B(n11076), .C(n2473), .D(n11290), .Q(n10677) );
  OAI222 U4270 ( .A(n2833), .B(n11074), .C(n2809), .D(n11289), .Q(n10684) );
  OAI222 U4273 ( .A(n2785), .B(n11072), .C(n2761), .D(n11288), .Q(n10683) );
  OAI222 U4276 ( .A(n2737), .B(n11070), .C(n2713), .D(n11287), .Q(n10682) );
  OAI222 U4279 ( .A(n2689), .B(n11068), .C(n2665), .D(n11286), .Q(n10681) );
  OAI222 U4284 ( .A(n3025), .B(n11066), .C(n3001), .D(n11285), .Q(n10691) );
  OAI222 U4287 ( .A(n2977), .B(n11064), .C(n2953), .D(n11284), .Q(n10690) );
  OAI222 U4290 ( .A(n2929), .B(n11062), .C(n2905), .D(n11283), .Q(n10689) );
  OAI222 U4293 ( .A(n2881), .B(n11060), .C(n2857), .D(n11282), .Q(n10688) );
  OAI222 U4298 ( .A(n1681), .B(n11058), .C(n1657), .D(n11281), .Q(n10699) );
  OAI222 U4301 ( .A(n1633), .B(n11056), .C(n1609), .D(n11280), .Q(n10698) );
  OAI222 U4304 ( .A(n1585), .B(n11054), .C(n1561), .D(n11279), .Q(n10697) );
  OAI222 U4307 ( .A(n1537), .B(n11052), .C(n1513), .D(n11278), .Q(n10696) );
  OAI222 U4311 ( .A(n1873), .B(n11050), .C(n1849), .D(n11277), .Q(n10703) );
  OAI222 U4314 ( .A(n1825), .B(n11048), .C(n1801), .D(n11276), .Q(n10702) );
  OAI222 U4317 ( .A(n1777), .B(n11046), .C(n1753), .D(n11275), .Q(n10701) );
  OAI222 U4320 ( .A(n1729), .B(n11044), .C(n1705), .D(n11274), .Q(n10700) );
  OAI222 U4324 ( .A(n2065), .B(n11042), .C(n2041), .D(n11273), .Q(n10707) );
  OAI222 U4327 ( .A(n2017), .B(n11040), .C(n1993), .D(n11272), .Q(n10706) );
  OAI222 U4330 ( .A(n1969), .B(n11038), .C(n1945), .D(n11271), .Q(n10705) );
  OAI222 U4333 ( .A(n1921), .B(n11036), .C(n1897), .D(n11270), .Q(n10704) );
  OAI222 U4338 ( .A(n2257), .B(n11034), .C(n2233), .D(n11269), .Q(n10713) );
  OAI222 U4341 ( .A(n2209), .B(n11032), .C(n2185), .D(n11268), .Q(n10712) );
  OAI222 U4344 ( .A(n2161), .B(n11030), .C(n2137), .D(n11267), .Q(n10711) );
  OAI222 U4347 ( .A(n2113), .B(n11028), .C(n2089), .D(n11266), .Q(n10710) );
  OAI222 U4353 ( .A(n913), .B(n11026), .C(n889), .D(n11265), .Q(n10723) );
  OAI222 U4356 ( .A(n865), .B(n11024), .C(n841), .D(n11264), .Q(n10722) );
  OAI222 U4359 ( .A(n817), .B(n11022), .C(n793), .D(n11263), .Q(n10721) );
  OAI222 U4362 ( .A(n769), .B(n11020), .C(n745), .D(n11262), .Q(n10720) );
  OAI222 U4366 ( .A(n1105), .B(n11018), .C(n1081), .D(n11261), .Q(n10727) );
  OAI222 U4369 ( .A(n1057), .B(n11016), .C(n1033), .D(n11260), .Q(n10726) );
  OAI222 U4372 ( .A(n1009), .B(n11014), .C(n985), .D(n11259), .Q(n10725) );
  OAI222 U4375 ( .A(n961), .B(n11012), .C(n937), .D(n11258), .Q(n10724) );
  OAI222 U4379 ( .A(n1297), .B(n11010), .C(n1273), .D(n11257), .Q(n10731) );
  OAI222 U4382 ( .A(n1249), .B(n11008), .C(n1225), .D(n11256), .Q(n10730) );
  OAI222 U4385 ( .A(n1201), .B(n11006), .C(n1177), .D(n11255), .Q(n10729) );
  OAI222 U4388 ( .A(n1153), .B(n11004), .C(n1129), .D(n11254), .Q(n10728) );
  OAI222 U4393 ( .A(n1489), .B(n11002), .C(n1465), .D(n11253), .Q(n10737) );
  OAI222 U4396 ( .A(n1441), .B(n11000), .C(n1417), .D(n11252), .Q(n10736) );
  OAI222 U4399 ( .A(n1393), .B(n10998), .C(n1369), .D(n11251), .Q(n10735) );
  OAI222 U4402 ( .A(n1345), .B(n10996), .C(n1321), .D(n11250), .Q(n10734) );
  OAI222 U4408 ( .A(n145), .B(n10994), .C(n121), .D(n11249), .Q(n10747) );
  OAI222 U4411 ( .A(n97), .B(n10992), .C(n73), .D(n11248), .Q(n10746) );
  OAI222 U4414 ( .A(n49), .B(n10990), .C(n25), .D(n11247), .Q(n10745) );
  OAI222 U4417 ( .A(n1), .B(n10988), .C(n6121), .D(n11246), .Q(n10744) );
  OAI222 U4421 ( .A(n337), .B(n10986), .C(n313), .D(n11245), .Q(n10751) );
  OAI222 U4424 ( .A(n289), .B(n10984), .C(n265), .D(n11244), .Q(n10750) );
  OAI222 U4427 ( .A(n241), .B(n10982), .C(n217), .D(n11243), .Q(n10749) );
  OAI222 U4430 ( .A(n193), .B(n10980), .C(n169), .D(n11242), .Q(n10748) );
  OAI222 U4434 ( .A(n529), .B(n10978), .C(n505), .D(n11241), .Q(n10755) );
  OAI222 U4437 ( .A(n481), .B(n10976), .C(n457), .D(n11240), .Q(n10754) );
  OAI222 U4440 ( .A(n433), .B(n10974), .C(n409), .D(n11239), .Q(n10753) );
  OAI222 U4443 ( .A(n385), .B(n10972), .C(n361), .D(n11238), .Q(n10752) );
  OAI222 U4448 ( .A(n721), .B(n10970), .C(n697), .D(n11237), .Q(n10760) );
  OAI222 U4451 ( .A(n673), .B(n10968), .C(n649), .D(n11236), .Q(n10759) );
  OAI222 U4454 ( .A(n625), .B(n10966), .C(n601), .D(n11235), .Q(n10758) );
  OAI222 U4457 ( .A(n577), .B(n10964), .C(n553), .D(n11234), .Q(n10757) );
  OAI222 U4465 ( .A(n5521), .B(n10962), .C(n5497), .D(n11233), .Q(n10773) );
  OAI222 U4468 ( .A(n5473), .B(n10960), .C(n5449), .D(n11232), .Q(n10772) );
  OAI222 U4471 ( .A(n5425), .B(n10958), .C(n5401), .D(n11231), .Q(n10771) );
  OAI222 U4474 ( .A(n5377), .B(n10956), .C(n5353), .D(n11230), .Q(n10770) );
  OAI222 U4478 ( .A(n5713), .B(n10954), .C(n5689), .D(n11229), .Q(n10777) );
  OAI222 U4481 ( .A(n5665), .B(n10952), .C(n5641), .D(n11228), .Q(n10776) );
  OAI222 U4484 ( .A(n5617), .B(n10950), .C(n5593), .D(n11227), .Q(n10775) );
  OAI222 U4487 ( .A(n5569), .B(n10948), .C(n5545), .D(n11226), .Q(n10774) );
  OAI222 U4491 ( .A(n5905), .B(n10946), .C(n5881), .D(n11225), .Q(n10781) );
  OAI222 U4494 ( .A(n5857), .B(n10944), .C(n5833), .D(n11224), .Q(n10780) );
  OAI222 U4497 ( .A(n5809), .B(n10942), .C(n5785), .D(n11223), .Q(n10779) );
  OAI222 U4500 ( .A(n5761), .B(n10940), .C(n5737), .D(n11222), .Q(n10778) );
  OAI222 U4505 ( .A(n6097), .B(n10938), .C(n6073), .D(n11221), .Q(n10787) );
  OAI222 U4508 ( .A(n6049), .B(n10936), .C(n6025), .D(n11220), .Q(n10786) );
  OAI222 U4511 ( .A(n6001), .B(n10934), .C(n5977), .D(n11219), .Q(n10785) );
  OAI222 U4514 ( .A(n5953), .B(n10932), .C(n5929), .D(n11218), .Q(n10784) );
  OAI222 U4520 ( .A(n4753), .B(n10930), .C(n4729), .D(n11217), .Q(n10796) );
  OAI222 U4523 ( .A(n4705), .B(n10928), .C(n4681), .D(n11216), .Q(n10795) );
  OAI222 U4526 ( .A(n4657), .B(n10926), .C(n4633), .D(n11215), .Q(n10794) );
  OAI222 U4529 ( .A(n4609), .B(n10924), .C(n4585), .D(n11214), .Q(n10793) );
  OAI222 U4533 ( .A(n4945), .B(n10922), .C(n4921), .D(n11213), .Q(n10800) );
  OAI222 U4536 ( .A(n4897), .B(n10920), .C(n4873), .D(n11212), .Q(n10799) );
  OAI222 U4539 ( .A(n4849), .B(n10918), .C(n4825), .D(n11211), .Q(n10798) );
  OAI222 U4542 ( .A(n4801), .B(n10916), .C(n4777), .D(n11210), .Q(n10797) );
  OAI222 U4546 ( .A(n5137), .B(n10914), .C(n5113), .D(n11209), .Q(n10804) );
  OAI222 U4549 ( .A(n5089), .B(n10912), .C(n5065), .D(n11208), .Q(n10803) );
  OAI222 U4552 ( .A(n5041), .B(n10910), .C(n5017), .D(n11207), .Q(n10802) );
  OAI222 U4555 ( .A(n4993), .B(n10908), .C(n4969), .D(n11206), .Q(n10801) );
  OAI222 U4560 ( .A(n5329), .B(n10906), .C(n5305), .D(n11205), .Q(n10809) );
  OAI222 U4563 ( .A(n5281), .B(n10904), .C(n5257), .D(n11204), .Q(n10808) );
  OAI222 U4566 ( .A(n5233), .B(n10902), .C(n5209), .D(n11203), .Q(n10807) );
  OAI222 U4569 ( .A(n5185), .B(n10900), .C(n5161), .D(n11202), .Q(n10806) );
  OAI222 U4576 ( .A(n3985), .B(n10898), .C(n3961), .D(n11201), .Q(n10818) );
  OAI222 U4579 ( .A(n3937), .B(n10896), .C(n3913), .D(n11200), .Q(n10817) );
  OAI222 U4582 ( .A(n3889), .B(n10894), .C(n3865), .D(n11199), .Q(n10816) );
  OAI222 U4585 ( .A(n3841), .B(n10892), .C(n3817), .D(n11198), .Q(n10815) );
  OAI222 U4589 ( .A(n4177), .B(n10890), .C(n4153), .D(n11197), .Q(n10822) );
  OAI222 U4592 ( .A(n4129), .B(n10888), .C(n4105), .D(n11196), .Q(n10821) );
  OAI222 U4595 ( .A(n4081), .B(n10886), .C(n4057), .D(n11195), .Q(n10820) );
  OAI222 U4598 ( .A(n4033), .B(n10884), .C(n4009), .D(n11194), .Q(n10819) );
  OAI222 U4602 ( .A(n4369), .B(n10882), .C(n4345), .D(n11193), .Q(n10826) );
  OAI222 U4605 ( .A(n4321), .B(n6192), .C(n4297), .D(n11192), .Q(n10825) );
  OAI222 U4608 ( .A(n4273), .B(n6190), .C(n4249), .D(n11191), .Q(n10824) );
  OAI222 U4611 ( .A(n4225), .B(n6188), .C(n4201), .D(n11190), .Q(n10823) );
  OAI222 U4617 ( .A(n4561), .B(n6186), .C(n4537), .D(n11189), .Q(n10832) );
  OAI222 U4620 ( .A(n4513), .B(n6184), .C(n4489), .D(n11188), .Q(n10831) );
  OAI222 U4623 ( .A(n4465), .B(n6182), .C(n4441), .D(n11187), .Q(n10830) );
  OAI222 U4626 ( .A(n4417), .B(n6180), .C(n4393), .D(n11186), .Q(n10829) );
  OAI222 U4632 ( .A(n3217), .B(n6178), .C(n3193), .D(n11185), .Q(n10841) );
  OAI222 U4635 ( .A(n3169), .B(n6176), .C(n3145), .D(n11184), .Q(n10840) );
  OAI222 U4638 ( .A(n3121), .B(n6174), .C(n3097), .D(n11183), .Q(n10839) );
  OAI222 U4641 ( .A(n3073), .B(n6172), .C(n3049), .D(n11182), .Q(n10838) );
  OAI222 U4648 ( .A(n3409), .B(n6170), .C(n3385), .D(n11181), .Q(n10846) );
  OAI222 U4651 ( .A(n3361), .B(n6168), .C(n3337), .D(n11180), .Q(n10845) );
  OAI222 U4654 ( .A(n3313), .B(n6166), .C(n3289), .D(n11179), .Q(n10844) );
  OAI222 U4657 ( .A(n3265), .B(n6164), .C(n3241), .D(n11178), .Q(n10843) );
  OAI222 U4661 ( .A(n3601), .B(n6162), .C(n3577), .D(n11177), .Q(n10850) );
  OAI222 U4666 ( .A(n3553), .B(n6160), .C(n3529), .D(n11176), .Q(n10849) );
  OAI222 U4671 ( .A(n3505), .B(n6158), .C(n3481), .D(n11175), .Q(n10848) );
  OAI222 U4676 ( .A(n3457), .B(n6156), .C(n3433), .D(n11174), .Q(n10847) );
  OAI222 U4685 ( .A(n3793), .B(n6154), .C(n3769), .D(n11173), .Q(n10870) );
  OAI222 U4690 ( .A(n3745), .B(n6152), .C(n3721), .D(n11172), .Q(n10869) );
  OAI222 U4696 ( .A(n3697), .B(n6150), .C(n3673), .D(n11171), .Q(n10868) );
  OAI222 U4703 ( .A(n3649), .B(n6148), .C(n3625), .D(n11170), .Q(n10867) );
  DF3 Q_reg_23 ( .D(N791), .C(n11303), .Q(Q_23) );
  DF3 Q_reg_22 ( .D(N792), .C(n11303), .Q(Q_22) );
  DF3 Q_reg_21 ( .D(N793), .C(n11303), .Q(Q_21) );
  DF3 Q_reg_20 ( .D(N794), .C(n11303), .Q(Q_20) );
  DF3 Q_reg_19 ( .D(N795), .C(n11302), .Q(Q_19) );
  DF3 Q_reg_18 ( .D(N796), .C(n11302), .Q(Q_18) );
  DF3 Q_reg_17 ( .D(N797), .C(n11302), .Q(Q_17) );
  DF3 Q_reg_16 ( .D(N798), .C(n11302), .Q(Q_16) );
  DF3 Q_reg_15 ( .D(N799), .C(n11301), .Q(Q_15) );
  DF3 Q_reg_14 ( .D(N800), .C(n11301), .Q(Q_14) );
  DF3 Q_reg_13 ( .D(N801), .C(n11301), .Q(Q_13) );
  DF3 Q_reg_12 ( .D(N802), .C(n11301), .Q(Q_12) );
  DF3 Q_reg_11 ( .D(N803), .C(n11300), .Q(Q_11) );
  DF3 Q_reg_10 ( .D(N804), .C(n11300), .Q(Q_10) );
  DF3 Q_reg_9 ( .D(N805), .C(n11300), .Q(Q_9) );
  DF3 Q_reg_8 ( .D(N806), .C(n11300), .Q(Q_8) );
  DF3 Q_reg_7 ( .D(N807), .C(n11299), .Q(Q_7) );
  DF3 Q_reg_6 ( .D(N808), .C(n11299), .Q(Q_6) );
  DF3 Q_reg_5 ( .D(N809), .C(n11299), .Q(Q_5) );
  DF3 Q_reg_4 ( .D(N810), .C(n11299), .Q(Q_4) );
  DF3 Q_reg_3 ( .D(N811), .C(n11298), .Q(Q_3) );
  DF3 Q_reg_2 ( .D(N812), .C(n11298), .Q(Q_2) );
  DF3 Q_reg_1 ( .D(N813), .C(n11298), .Q(Q_1) );
  DF3 Q_reg_0 ( .D(N814), .C(n11298), .Q(Q_0) );
  DFE1 \mem_reg_15][23  ( .D(D_23), .E(n6437), .C(wclk), .QN(n5761) );
  DFE1 \mem_reg_15][22  ( .D(D_22), .E(n6437), .C(wclk), .QN(n5762) );
  DFE1 \mem_reg_15][21  ( .D(D_21), .E(n6437), .C(wclk), .QN(n5763) );
  DFE1 \mem_reg_15][20  ( .D(D_20), .E(n6437), .C(wclk), .QN(n5764) );
  DFE1 \mem_reg_15][19  ( .D(D_19), .E(n6437), .C(wclk), .QN(n5765) );
  DFE1 \mem_reg_15][18  ( .D(D_18), .E(n6437), .C(wclk), .QN(n5766) );
  DFE1 \mem_reg_15][17  ( .D(D_17), .E(n6437), .C(wclk), .QN(n5767) );
  DFE1 \mem_reg_15][16  ( .D(D_16), .E(n6437), .C(wclk), .QN(n5768) );
  DFE1 \mem_reg_15][15  ( .D(D_15), .E(n6437), .C(wclk), .QN(n5769) );
  DFE1 \mem_reg_15][14  ( .D(D_14), .E(n6437), .C(wclk), .QN(n5770) );
  DFE1 \mem_reg_15][13  ( .D(D_13), .E(n6437), .C(wclk), .QN(n5771) );
  DFE1 \mem_reg_15][12  ( .D(D_12), .E(n6437), .C(wclk), .QN(n5772) );
  DFE1 \mem_reg_15][11  ( .D(D_11), .E(n6437), .C(wclk), .QN(n5773) );
  DFE1 \mem_reg_15][10  ( .D(D_10), .E(n6437), .C(wclk), .QN(n5774) );
  DFE1 \mem_reg_15][9  ( .D(D_9), .E(n6437), .C(wclk), .QN(n5775) );
  DFE1 \mem_reg_15][8  ( .D(D_8), .E(n6437), .C(wclk), .QN(n5776) );
  DFE1 \mem_reg_15][7  ( .D(D_7), .E(n6437), .C(wclk), .QN(n5777) );
  DFE1 \mem_reg_15][6  ( .D(D_6), .E(n6437), .C(wclk), .QN(n5778) );
  DFE1 \mem_reg_15][5  ( .D(D_5), .E(n6437), .C(wclk), .QN(n5779) );
  DFE1 \mem_reg_15][4  ( .D(D_4), .E(n6437), .C(wclk), .QN(n5780) );
  DFE1 \mem_reg_15][3  ( .D(D_3), .E(n6437), .C(wclk), .QN(n5781) );
  DFE1 \mem_reg_15][2  ( .D(D_2), .E(n6437), .C(wclk), .QN(n5782) );
  DFE1 \mem_reg_15][1  ( .D(D_1), .E(n6437), .C(wclk), .QN(n5783) );
  DFE1 \mem_reg_15][0  ( .D(D_0), .E(n6437), .C(wclk), .QN(n5784) );
  DFE1 \mem_reg_14][23  ( .D(D_23), .E(n6436), .C(wclk), .QN(n5785) );
  DFE1 \mem_reg_14][22  ( .D(D_22), .E(n6436), .C(wclk), .QN(n5786) );
  DFE1 \mem_reg_14][21  ( .D(D_21), .E(n6436), .C(wclk), .QN(n5787) );
  DFE1 \mem_reg_14][20  ( .D(D_20), .E(n6436), .C(wclk), .QN(n5788) );
  DFE1 \mem_reg_14][19  ( .D(D_19), .E(n6436), .C(wclk), .QN(n5789) );
  DFE1 \mem_reg_14][18  ( .D(D_18), .E(n6436), .C(wclk), .QN(n5790) );
  DFE1 \mem_reg_14][17  ( .D(D_17), .E(n6436), .C(wclk), .QN(n5791) );
  DFE1 \mem_reg_14][16  ( .D(D_16), .E(n6436), .C(wclk), .QN(n5792) );
  DFE1 \mem_reg_14][15  ( .D(D_15), .E(n6436), .C(wclk), .QN(n5793) );
  DFE1 \mem_reg_14][14  ( .D(D_14), .E(n6436), .C(wclk), .QN(n5794) );
  DFE1 \mem_reg_14][13  ( .D(D_13), .E(n6436), .C(wclk), .QN(n5795) );
  DFE1 \mem_reg_14][12  ( .D(D_12), .E(n6436), .C(wclk), .QN(n5796) );
  DFE1 \mem_reg_14][11  ( .D(D_11), .E(n6436), .C(wclk), .QN(n5797) );
  DFE1 \mem_reg_14][10  ( .D(D_10), .E(n6436), .C(wclk), .QN(n5798) );
  DFE1 \mem_reg_14][9  ( .D(D_9), .E(n6436), .C(wclk), .QN(n5799) );
  DFE1 \mem_reg_14][8  ( .D(D_8), .E(n6436), .C(wclk), .QN(n5800) );
  DFE1 \mem_reg_14][7  ( .D(D_7), .E(n6436), .C(wclk), .QN(n5801) );
  DFE1 \mem_reg_14][6  ( .D(D_6), .E(n6436), .C(wclk), .QN(n5802) );
  DFE1 \mem_reg_14][5  ( .D(D_5), .E(n6436), .C(wclk), .QN(n5803) );
  DFE1 \mem_reg_14][4  ( .D(D_4), .E(n6436), .C(wclk), .QN(n5804) );
  DFE1 \mem_reg_14][3  ( .D(D_3), .E(n6436), .C(wclk), .QN(n5805) );
  DFE1 \mem_reg_14][2  ( .D(D_2), .E(n6436), .C(wclk), .QN(n5806) );
  DFE1 \mem_reg_14][1  ( .D(D_1), .E(n6436), .C(wclk), .QN(n5807) );
  DFE1 \mem_reg_14][0  ( .D(D_0), .E(n6436), .C(wclk), .QN(n5808) );
  DFE1 \mem_reg_12][23  ( .D(D_23), .E(n6433), .C(wclk), .QN(n5833) );
  DFE1 \mem_reg_12][22  ( .D(D_22), .E(n6433), .C(wclk), .QN(n5834) );
  DFE1 \mem_reg_12][21  ( .D(D_21), .E(n6433), .C(wclk), .QN(n5835) );
  DFE1 \mem_reg_12][20  ( .D(D_20), .E(n6433), .C(wclk), .QN(n5836) );
  DFE1 \mem_reg_12][19  ( .D(D_19), .E(n6433), .C(wclk), .QN(n5837) );
  DFE1 \mem_reg_12][18  ( .D(D_18), .E(n6433), .C(wclk), .QN(n5838) );
  DFE1 \mem_reg_12][17  ( .D(D_17), .E(n6433), .C(wclk), .QN(n5839) );
  DFE1 \mem_reg_12][16  ( .D(D_16), .E(n6433), .C(wclk), .QN(n5840) );
  DFE1 \mem_reg_12][15  ( .D(D_15), .E(n6433), .C(wclk), .QN(n5841) );
  DFE1 \mem_reg_12][14  ( .D(D_14), .E(n6433), .C(wclk), .QN(n5842) );
  DFE1 \mem_reg_12][13  ( .D(D_13), .E(n6433), .C(wclk), .QN(n5843) );
  DFE1 \mem_reg_12][12  ( .D(D_12), .E(n6433), .C(wclk), .QN(n5844) );
  DFE1 \mem_reg_12][11  ( .D(D_11), .E(n6433), .C(wclk), .QN(n5845) );
  DFE1 \mem_reg_12][10  ( .D(D_10), .E(n6433), .C(wclk), .QN(n5846) );
  DFE1 \mem_reg_12][9  ( .D(D_9), .E(n6433), .C(wclk), .QN(n5847) );
  DFE1 \mem_reg_12][8  ( .D(D_8), .E(n6433), .C(wclk), .QN(n5848) );
  DFE1 \mem_reg_12][7  ( .D(D_7), .E(n6433), .C(wclk), .QN(n5849) );
  DFE1 \mem_reg_12][6  ( .D(D_6), .E(n6433), .C(wclk), .QN(n5850) );
  DFE1 \mem_reg_12][5  ( .D(D_5), .E(n6433), .C(wclk), .QN(n5851) );
  DFE1 \mem_reg_12][4  ( .D(D_4), .E(n6433), .C(wclk), .QN(n5852) );
  DFE1 \mem_reg_12][3  ( .D(D_3), .E(n6433), .C(wclk), .QN(n5853) );
  DFE1 \mem_reg_12][2  ( .D(D_2), .E(n6433), .C(wclk), .QN(n5854) );
  DFE1 \mem_reg_12][1  ( .D(D_1), .E(n6433), .C(wclk), .QN(n5855) );
  DFE1 \mem_reg_12][0  ( .D(D_0), .E(n6433), .C(wclk), .QN(n5856) );
  DFE1 \mem_reg_9][23  ( .D(D_23), .E(n6430), .C(wclk), .QN(n5905) );
  DFE1 \mem_reg_9][22  ( .D(D_22), .E(n6430), .C(wclk), .QN(n5906) );
  DFE1 \mem_reg_9][21  ( .D(D_21), .E(n6430), .C(wclk), .QN(n5907) );
  DFE1 \mem_reg_9][20  ( .D(D_20), .E(n6430), .C(wclk), .QN(n5908) );
  DFE1 \mem_reg_9][19  ( .D(D_19), .E(n6430), .C(wclk), .QN(n5909) );
  DFE1 \mem_reg_9][18  ( .D(D_18), .E(n6430), .C(wclk), .QN(n5910) );
  DFE1 \mem_reg_9][17  ( .D(D_17), .E(n6430), .C(wclk), .QN(n5911) );
  DFE1 \mem_reg_9][16  ( .D(D_16), .E(n6430), .C(wclk), .QN(n5912) );
  DFE1 \mem_reg_9][15  ( .D(D_15), .E(n6430), .C(wclk), .QN(n5913) );
  DFE1 \mem_reg_9][14  ( .D(D_14), .E(n6430), .C(wclk), .QN(n5914) );
  DFE1 \mem_reg_9][13  ( .D(D_13), .E(n6430), .C(wclk), .QN(n5915) );
  DFE1 \mem_reg_9][12  ( .D(D_12), .E(n6430), .C(wclk), .QN(n5916) );
  DFE1 \mem_reg_9][11  ( .D(D_11), .E(n6430), .C(wclk), .QN(n5917) );
  DFE1 \mem_reg_9][10  ( .D(D_10), .E(n6430), .C(wclk), .QN(n5918) );
  DFE1 \mem_reg_9][9  ( .D(D_9), .E(n6430), .C(wclk), .QN(n5919) );
  DFE1 \mem_reg_9][8  ( .D(D_8), .E(n6430), .C(wclk), .QN(n5920) );
  DFE1 \mem_reg_9][7  ( .D(D_7), .E(n6430), .C(wclk), .QN(n5921) );
  DFE1 \mem_reg_9][6  ( .D(D_6), .E(n6430), .C(wclk), .QN(n5922) );
  DFE1 \mem_reg_9][5  ( .D(D_5), .E(n6430), .C(wclk), .QN(n5923) );
  DFE1 \mem_reg_9][4  ( .D(D_4), .E(n6430), .C(wclk), .QN(n5924) );
  DFE1 \mem_reg_9][3  ( .D(D_3), .E(n6430), .C(wclk), .QN(n5925) );
  DFE1 \mem_reg_9][2  ( .D(D_2), .E(n6430), .C(wclk), .QN(n5926) );
  DFE1 \mem_reg_9][1  ( .D(D_1), .E(n6430), .C(wclk), .QN(n5927) );
  DFE1 \mem_reg_9][0  ( .D(D_0), .E(n6430), .C(wclk), .QN(n5928) );
  DFE1 \mem_reg_8][23  ( .D(D_23), .E(n6429), .C(wclk), .QN(n5929) );
  DFE1 \mem_reg_8][22  ( .D(D_22), .E(n6429), .C(wclk), .QN(n5930) );
  DFE1 \mem_reg_8][21  ( .D(D_21), .E(n6429), .C(wclk), .QN(n5931) );
  DFE1 \mem_reg_8][20  ( .D(D_20), .E(n6429), .C(wclk), .QN(n5932) );
  DFE1 \mem_reg_8][19  ( .D(D_19), .E(n6429), .C(wclk), .QN(n5933) );
  DFE1 \mem_reg_8][18  ( .D(D_18), .E(n6429), .C(wclk), .QN(n5934) );
  DFE1 \mem_reg_8][17  ( .D(D_17), .E(n6429), .C(wclk), .QN(n5935) );
  DFE1 \mem_reg_8][16  ( .D(D_16), .E(n6429), .C(wclk), .QN(n5936) );
  DFE1 \mem_reg_8][15  ( .D(D_15), .E(n6429), .C(wclk), .QN(n5937) );
  DFE1 \mem_reg_8][14  ( .D(D_14), .E(n6429), .C(wclk), .QN(n5938) );
  DFE1 \mem_reg_8][13  ( .D(D_13), .E(n6429), .C(wclk), .QN(n5939) );
  DFE1 \mem_reg_8][12  ( .D(D_12), .E(n6429), .C(wclk), .QN(n5940) );
  DFE1 \mem_reg_8][11  ( .D(D_11), .E(n6429), .C(wclk), .QN(n5941) );
  DFE1 \mem_reg_8][10  ( .D(D_10), .E(n6429), .C(wclk), .QN(n5942) );
  DFE1 \mem_reg_8][9  ( .D(D_9), .E(n6429), .C(wclk), .QN(n5943) );
  DFE1 \mem_reg_8][8  ( .D(D_8), .E(n6429), .C(wclk), .QN(n5944) );
  DFE1 \mem_reg_8][7  ( .D(D_7), .E(n6429), .C(wclk), .QN(n5945) );
  DFE1 \mem_reg_8][6  ( .D(D_6), .E(n6429), .C(wclk), .QN(n5946) );
  DFE1 \mem_reg_8][5  ( .D(D_5), .E(n6429), .C(wclk), .QN(n5947) );
  DFE1 \mem_reg_8][4  ( .D(D_4), .E(n6429), .C(wclk), .QN(n5948) );
  DFE1 \mem_reg_8][3  ( .D(D_3), .E(n6429), .C(wclk), .QN(n5949) );
  DFE1 \mem_reg_8][2  ( .D(D_2), .E(n6429), .C(wclk), .QN(n5950) );
  DFE1 \mem_reg_8][1  ( .D(D_1), .E(n6429), .C(wclk), .QN(n5951) );
  DFE1 \mem_reg_8][0  ( .D(D_0), .E(n6429), .C(wclk), .QN(n5952) );
  DFE1 \mem_reg_7][23  ( .D(D_23), .E(n6428), .C(wclk), .QN(n5953) );
  DFE1 \mem_reg_7][22  ( .D(D_22), .E(n6428), .C(wclk), .QN(n5954) );
  DFE1 \mem_reg_7][21  ( .D(D_21), .E(n6428), .C(wclk), .QN(n5955) );
  DFE1 \mem_reg_7][20  ( .D(D_20), .E(n6428), .C(wclk), .QN(n5956) );
  DFE1 \mem_reg_7][19  ( .D(D_19), .E(n6428), .C(wclk), .QN(n5957) );
  DFE1 \mem_reg_7][18  ( .D(D_18), .E(n6428), .C(wclk), .QN(n5958) );
  DFE1 \mem_reg_7][17  ( .D(D_17), .E(n6428), .C(wclk), .QN(n5959) );
  DFE1 \mem_reg_7][16  ( .D(D_16), .E(n6428), .C(wclk), .QN(n5960) );
  DFE1 \mem_reg_7][15  ( .D(D_15), .E(n6428), .C(wclk), .QN(n5961) );
  DFE1 \mem_reg_7][14  ( .D(D_14), .E(n6428), .C(wclk), .QN(n5962) );
  DFE1 \mem_reg_7][13  ( .D(D_13), .E(n6428), .C(wclk), .QN(n5963) );
  DFE1 \mem_reg_7][12  ( .D(D_12), .E(n6428), .C(wclk), .QN(n5964) );
  DFE1 \mem_reg_7][11  ( .D(D_11), .E(n6428), .C(wclk), .QN(n5965) );
  DFE1 \mem_reg_7][10  ( .D(D_10), .E(n6428), .C(wclk), .QN(n5966) );
  DFE1 \mem_reg_7][9  ( .D(D_9), .E(n6428), .C(wclk), .QN(n5967) );
  DFE1 \mem_reg_7][8  ( .D(D_8), .E(n6428), .C(wclk), .QN(n5968) );
  DFE1 \mem_reg_7][7  ( .D(D_7), .E(n6428), .C(wclk), .QN(n5969) );
  DFE1 \mem_reg_7][6  ( .D(D_6), .E(n6428), .C(wclk), .QN(n5970) );
  DFE1 \mem_reg_7][5  ( .D(D_5), .E(n6428), .C(wclk), .QN(n5971) );
  DFE1 \mem_reg_7][4  ( .D(D_4), .E(n6428), .C(wclk), .QN(n5972) );
  DFE1 \mem_reg_7][3  ( .D(D_3), .E(n6428), .C(wclk), .QN(n5973) );
  DFE1 \mem_reg_7][2  ( .D(D_2), .E(n6428), .C(wclk), .QN(n5974) );
  DFE1 \mem_reg_7][1  ( .D(D_1), .E(n6428), .C(wclk), .QN(n5975) );
  DFE1 \mem_reg_7][0  ( .D(D_0), .E(n6428), .C(wclk), .QN(n5976) );
  DFE1 \mem_reg_6][23  ( .D(D_23), .E(n6427), .C(wclk), .QN(n5977) );
  DFE1 \mem_reg_6][22  ( .D(D_22), .E(n6427), .C(wclk), .QN(n5978) );
  DFE1 \mem_reg_6][21  ( .D(D_21), .E(n6427), .C(wclk), .QN(n5979) );
  DFE1 \mem_reg_6][20  ( .D(D_20), .E(n6427), .C(wclk), .QN(n5980) );
  DFE1 \mem_reg_6][19  ( .D(D_19), .E(n6427), .C(wclk), .QN(n5981) );
  DFE1 \mem_reg_6][18  ( .D(D_18), .E(n6427), .C(wclk), .QN(n5982) );
  DFE1 \mem_reg_6][17  ( .D(D_17), .E(n6427), .C(wclk), .QN(n5983) );
  DFE1 \mem_reg_6][16  ( .D(D_16), .E(n6427), .C(wclk), .QN(n5984) );
  DFE1 \mem_reg_6][15  ( .D(D_15), .E(n6427), .C(wclk), .QN(n5985) );
  DFE1 \mem_reg_6][14  ( .D(D_14), .E(n6427), .C(wclk), .QN(n5986) );
  DFE1 \mem_reg_6][13  ( .D(D_13), .E(n6427), .C(wclk), .QN(n5987) );
  DFE1 \mem_reg_6][12  ( .D(D_12), .E(n6427), .C(wclk), .QN(n5988) );
  DFE1 \mem_reg_6][11  ( .D(D_11), .E(n6427), .C(wclk), .QN(n5989) );
  DFE1 \mem_reg_6][10  ( .D(D_10), .E(n6427), .C(wclk), .QN(n5990) );
  DFE1 \mem_reg_6][9  ( .D(D_9), .E(n6427), .C(wclk), .QN(n5991) );
  DFE1 \mem_reg_6][8  ( .D(D_8), .E(n6427), .C(wclk), .QN(n5992) );
  DFE1 \mem_reg_6][7  ( .D(D_7), .E(n6427), .C(wclk), .QN(n5993) );
  DFE1 \mem_reg_6][6  ( .D(D_6), .E(n6427), .C(wclk), .QN(n5994) );
  DFE1 \mem_reg_6][5  ( .D(D_5), .E(n6427), .C(wclk), .QN(n5995) );
  DFE1 \mem_reg_6][4  ( .D(D_4), .E(n6427), .C(wclk), .QN(n5996) );
  DFE1 \mem_reg_6][3  ( .D(D_3), .E(n6427), .C(wclk), .QN(n5997) );
  DFE1 \mem_reg_6][2  ( .D(D_2), .E(n6427), .C(wclk), .QN(n5998) );
  DFE1 \mem_reg_6][1  ( .D(D_1), .E(n6427), .C(wclk), .QN(n5999) );
  DFE1 \mem_reg_6][0  ( .D(D_0), .E(n6427), .C(wclk), .QN(n6000) );
  DFE1 \mem_reg_4][23  ( .D(D_23), .E(n6425), .C(wclk), .QN(n6025) );
  DFE1 \mem_reg_4][22  ( .D(D_22), .E(n6425), .C(wclk), .QN(n6026) );
  DFE1 \mem_reg_4][21  ( .D(D_21), .E(n6425), .C(wclk), .QN(n6027) );
  DFE1 \mem_reg_4][20  ( .D(D_20), .E(n6425), .C(wclk), .QN(n6028) );
  DFE1 \mem_reg_4][19  ( .D(D_19), .E(n6425), .C(wclk), .QN(n6029) );
  DFE1 \mem_reg_4][18  ( .D(D_18), .E(n6425), .C(wclk), .QN(n6030) );
  DFE1 \mem_reg_4][17  ( .D(D_17), .E(n6425), .C(wclk), .QN(n6031) );
  DFE1 \mem_reg_4][16  ( .D(D_16), .E(n6425), .C(wclk), .QN(n6032) );
  DFE1 \mem_reg_4][15  ( .D(D_15), .E(n6425), .C(wclk), .QN(n6033) );
  DFE1 \mem_reg_4][14  ( .D(D_14), .E(n6425), .C(wclk), .QN(n6034) );
  DFE1 \mem_reg_4][13  ( .D(D_13), .E(n6425), .C(wclk), .QN(n6035) );
  DFE1 \mem_reg_4][12  ( .D(D_12), .E(n6425), .C(wclk), .QN(n6036) );
  DFE1 \mem_reg_4][11  ( .D(D_11), .E(n6425), .C(wclk), .QN(n6037) );
  DFE1 \mem_reg_4][10  ( .D(D_10), .E(n6425), .C(wclk), .QN(n6038) );
  DFE1 \mem_reg_4][9  ( .D(D_9), .E(n6425), .C(wclk), .QN(n6039) );
  DFE1 \mem_reg_4][8  ( .D(D_8), .E(n6425), .C(wclk), .QN(n6040) );
  DFE1 \mem_reg_4][7  ( .D(D_7), .E(n6425), .C(wclk), .QN(n6041) );
  DFE1 \mem_reg_4][6  ( .D(D_6), .E(n6425), .C(wclk), .QN(n6042) );
  DFE1 \mem_reg_4][5  ( .D(D_5), .E(n6425), .C(wclk), .QN(n6043) );
  DFE1 \mem_reg_4][4  ( .D(D_4), .E(n6425), .C(wclk), .QN(n6044) );
  DFE1 \mem_reg_4][3  ( .D(D_3), .E(n6425), .C(wclk), .QN(n6045) );
  DFE1 \mem_reg_4][2  ( .D(D_2), .E(n6425), .C(wclk), .QN(n6046) );
  DFE1 \mem_reg_4][1  ( .D(D_1), .E(n6425), .C(wclk), .QN(n6047) );
  DFE1 \mem_reg_4][0  ( .D(D_0), .E(n6425), .C(wclk), .QN(n6048) );
  DFE1 \mem_reg_3][23  ( .D(D_23), .E(n6423), .C(wclk), .QN(n6049) );
  DFE1 \mem_reg_3][22  ( .D(D_22), .E(n6423), .C(wclk), .QN(n6050) );
  DFE1 \mem_reg_3][21  ( .D(D_21), .E(n6423), .C(wclk), .QN(n6051) );
  DFE1 \mem_reg_3][20  ( .D(D_20), .E(n6423), .C(wclk), .QN(n6052) );
  DFE1 \mem_reg_3][19  ( .D(D_19), .E(n6423), .C(wclk), .QN(n6053) );
  DFE1 \mem_reg_3][18  ( .D(D_18), .E(n6423), .C(wclk), .QN(n6054) );
  DFE1 \mem_reg_3][17  ( .D(D_17), .E(n6423), .C(wclk), .QN(n6055) );
  DFE1 \mem_reg_3][16  ( .D(D_16), .E(n6423), .C(wclk), .QN(n6056) );
  DFE1 \mem_reg_3][15  ( .D(D_15), .E(n6423), .C(wclk), .QN(n6057) );
  DFE1 \mem_reg_3][14  ( .D(D_14), .E(n6423), .C(wclk), .QN(n6058) );
  DFE1 \mem_reg_3][13  ( .D(D_13), .E(n6423), .C(wclk), .QN(n6059) );
  DFE1 \mem_reg_3][12  ( .D(D_12), .E(n6423), .C(wclk), .QN(n6060) );
  DFE1 \mem_reg_3][11  ( .D(D_11), .E(n6423), .C(wclk), .QN(n6061) );
  DFE1 \mem_reg_3][10  ( .D(D_10), .E(n6423), .C(wclk), .QN(n6062) );
  DFE1 \mem_reg_3][9  ( .D(D_9), .E(n6423), .C(wclk), .QN(n6063) );
  DFE1 \mem_reg_3][8  ( .D(D_8), .E(n6423), .C(wclk), .QN(n6064) );
  DFE1 \mem_reg_3][7  ( .D(D_7), .E(n6423), .C(wclk), .QN(n6065) );
  DFE1 \mem_reg_3][6  ( .D(D_6), .E(n6423), .C(wclk), .QN(n6066) );
  DFE1 \mem_reg_3][5  ( .D(D_5), .E(n6423), .C(wclk), .QN(n6067) );
  DFE1 \mem_reg_3][4  ( .D(D_4), .E(n6423), .C(wclk), .QN(n6068) );
  DFE1 \mem_reg_3][3  ( .D(D_3), .E(n6423), .C(wclk), .QN(n6069) );
  DFE1 \mem_reg_3][2  ( .D(D_2), .E(n6423), .C(wclk), .QN(n6070) );
  DFE1 \mem_reg_3][1  ( .D(D_1), .E(n6423), .C(wclk), .QN(n6071) );
  DFE1 \mem_reg_3][0  ( .D(D_0), .E(n6423), .C(wclk), .QN(n6072) );
  DFE1 \mem_reg_2][23  ( .D(D_23), .E(n6422), .C(wclk), .QN(n6073) );
  DFE1 \mem_reg_2][22  ( .D(D_22), .E(n6422), .C(wclk), .QN(n6074) );
  DFE1 \mem_reg_2][21  ( .D(D_21), .E(n6422), .C(wclk), .QN(n6075) );
  DFE1 \mem_reg_2][20  ( .D(D_20), .E(n6422), .C(wclk), .QN(n6076) );
  DFE1 \mem_reg_2][19  ( .D(D_19), .E(n6422), .C(wclk), .QN(n6077) );
  DFE1 \mem_reg_2][18  ( .D(D_18), .E(n6422), .C(wclk), .QN(n6078) );
  DFE1 \mem_reg_2][17  ( .D(D_17), .E(n6422), .C(wclk), .QN(n6079) );
  DFE1 \mem_reg_2][16  ( .D(D_16), .E(n6422), .C(wclk), .QN(n6080) );
  DFE1 \mem_reg_2][15  ( .D(D_15), .E(n6422), .C(wclk), .QN(n6081) );
  DFE1 \mem_reg_2][14  ( .D(D_14), .E(n6422), .C(wclk), .QN(n6082) );
  DFE1 \mem_reg_2][13  ( .D(D_13), .E(n6422), .C(wclk), .QN(n6083) );
  DFE1 \mem_reg_2][12  ( .D(D_12), .E(n6422), .C(wclk), .QN(n6084) );
  DFE1 \mem_reg_2][11  ( .D(D_11), .E(n6422), .C(wclk), .QN(n6085) );
  DFE1 \mem_reg_2][10  ( .D(D_10), .E(n6422), .C(wclk), .QN(n6086) );
  DFE1 \mem_reg_2][9  ( .D(D_9), .E(n6422), .C(wclk), .QN(n6087) );
  DFE1 \mem_reg_2][8  ( .D(D_8), .E(n6422), .C(wclk), .QN(n6088) );
  DFE1 \mem_reg_2][7  ( .D(D_7), .E(n6422), .C(wclk), .QN(n6089) );
  DFE1 \mem_reg_2][6  ( .D(D_6), .E(n6422), .C(wclk), .QN(n6090) );
  DFE1 \mem_reg_2][5  ( .D(D_5), .E(n6422), .C(wclk), .QN(n6091) );
  DFE1 \mem_reg_2][4  ( .D(D_4), .E(n6422), .C(wclk), .QN(n6092) );
  DFE1 \mem_reg_2][3  ( .D(D_3), .E(n6422), .C(wclk), .QN(n6093) );
  DFE1 \mem_reg_2][2  ( .D(D_2), .E(n6422), .C(wclk), .QN(n6094) );
  DFE1 \mem_reg_2][1  ( .D(D_1), .E(n6422), .C(wclk), .QN(n6095) );
  DFE1 \mem_reg_2][0  ( .D(D_0), .E(n6422), .C(wclk), .QN(n6096) );
  DFE1 \mem_reg_0][23  ( .D(D_23), .E(n6419), .C(wclk), .QN(n6121) );
  DFE1 \mem_reg_0][22  ( .D(D_22), .E(n6419), .C(wclk), .QN(n6122) );
  DFE1 \mem_reg_0][21  ( .D(D_21), .E(n6419), .C(wclk), .QN(n6123) );
  DFE1 \mem_reg_0][20  ( .D(D_20), .E(n6419), .C(wclk), .QN(n6124) );
  DFE1 \mem_reg_0][19  ( .D(D_19), .E(n6419), .C(wclk), .QN(n6125) );
  DFE1 \mem_reg_0][18  ( .D(D_18), .E(n6419), .C(wclk), .QN(n6126) );
  DFE1 \mem_reg_0][17  ( .D(D_17), .E(n6419), .C(wclk), .QN(n6127) );
  DFE1 \mem_reg_0][16  ( .D(D_16), .E(n6419), .C(wclk), .QN(n6128) );
  DFE1 \mem_reg_0][15  ( .D(D_15), .E(n6419), .C(wclk), .QN(n6129) );
  DFE1 \mem_reg_0][14  ( .D(D_14), .E(n6419), .C(wclk), .QN(n6130) );
  DFE1 \mem_reg_0][13  ( .D(D_13), .E(n6419), .C(wclk), .QN(n6131) );
  DFE1 \mem_reg_0][12  ( .D(D_12), .E(n6419), .C(wclk), .QN(n6132) );
  DFE1 \mem_reg_0][11  ( .D(D_11), .E(n6419), .C(wclk), .QN(n6133) );
  DFE1 \mem_reg_0][10  ( .D(D_10), .E(n6419), .C(wclk), .QN(n6134) );
  DFE1 \mem_reg_0][9  ( .D(D_9), .E(n6419), .C(wclk), .QN(n6135) );
  DFE1 \mem_reg_0][8  ( .D(D_8), .E(n6419), .C(wclk), .QN(n6136) );
  DFE1 \mem_reg_0][7  ( .D(D_7), .E(n6419), .C(wclk), .QN(n6137) );
  DFE1 \mem_reg_0][6  ( .D(D_6), .E(n6419), .C(wclk), .QN(n6138) );
  DFE1 \mem_reg_0][5  ( .D(D_5), .E(n6419), .C(wclk), .QN(n6139) );
  DFE1 \mem_reg_0][4  ( .D(D_4), .E(n6419), .C(wclk), .QN(n6140) );
  DFE1 \mem_reg_0][3  ( .D(D_3), .E(n6419), .C(wclk), .QN(n6141) );
  DFE1 \mem_reg_0][2  ( .D(D_2), .E(n6419), .C(wclk), .QN(n6142) );
  DFE1 \mem_reg_0][1  ( .D(D_1), .E(n6419), .C(wclk), .QN(n6143) );
  DFE1 \mem_reg_0][0  ( .D(D_0), .E(n6419), .C(wclk), .QN(n6144) );
  DFE1 \mem_reg_11][23  ( .D(D_23), .E(n6432), .C(wclk), .QN(n5857) );
  DFE1 \mem_reg_11][22  ( .D(D_22), .E(n6432), .C(wclk), .QN(n5858) );
  DFE1 \mem_reg_11][21  ( .D(D_21), .E(n6432), .C(wclk), .QN(n5859) );
  DFE1 \mem_reg_11][20  ( .D(D_20), .E(n6432), .C(wclk), .QN(n5860) );
  DFE1 \mem_reg_11][19  ( .D(D_19), .E(n6432), .C(wclk), .QN(n5861) );
  DFE1 \mem_reg_11][18  ( .D(D_18), .E(n6432), .C(wclk), .QN(n5862) );
  DFE1 \mem_reg_11][17  ( .D(D_17), .E(n6432), .C(wclk), .QN(n5863) );
  DFE1 \mem_reg_11][16  ( .D(D_16), .E(n6432), .C(wclk), .QN(n5864) );
  DFE1 \mem_reg_11][15  ( .D(D_15), .E(n6432), .C(wclk), .QN(n5865) );
  DFE1 \mem_reg_11][14  ( .D(D_14), .E(n6432), .C(wclk), .QN(n5866) );
  DFE1 \mem_reg_11][13  ( .D(D_13), .E(n6432), .C(wclk), .QN(n5867) );
  DFE1 \mem_reg_11][12  ( .D(D_12), .E(n6432), .C(wclk), .QN(n5868) );
  DFE1 \mem_reg_11][11  ( .D(D_11), .E(n6432), .C(wclk), .QN(n5869) );
  DFE1 \mem_reg_11][10  ( .D(D_10), .E(n6432), .C(wclk), .QN(n5870) );
  DFE1 \mem_reg_11][9  ( .D(D_9), .E(n6432), .C(wclk), .QN(n5871) );
  DFE1 \mem_reg_11][8  ( .D(D_8), .E(n6432), .C(wclk), .QN(n5872) );
  DFE1 \mem_reg_11][7  ( .D(D_7), .E(n6432), .C(wclk), .QN(n5873) );
  DFE1 \mem_reg_11][6  ( .D(D_6), .E(n6432), .C(wclk), .QN(n5874) );
  DFE1 \mem_reg_11][5  ( .D(D_5), .E(n6432), .C(wclk), .QN(n5875) );
  DFE1 \mem_reg_11][4  ( .D(D_4), .E(n6432), .C(wclk), .QN(n5876) );
  DFE1 \mem_reg_11][3  ( .D(D_3), .E(n6432), .C(wclk), .QN(n5877) );
  DFE1 \mem_reg_11][2  ( .D(D_2), .E(n6432), .C(wclk), .QN(n5878) );
  DFE1 \mem_reg_11][1  ( .D(D_1), .E(n6432), .C(wclk), .QN(n5879) );
  DFE1 \mem_reg_11][0  ( .D(D_0), .E(n6432), .C(wclk), .QN(n5880) );
  DFE1 \mem_reg_10][23  ( .D(D_23), .E(n6431), .C(wclk), .QN(n5881) );
  DFE1 \mem_reg_10][22  ( .D(D_22), .E(n6431), .C(wclk), .QN(n5882) );
  DFE1 \mem_reg_10][21  ( .D(D_21), .E(n6431), .C(wclk), .QN(n5883) );
  DFE1 \mem_reg_10][20  ( .D(D_20), .E(n6431), .C(wclk), .QN(n5884) );
  DFE1 \mem_reg_10][19  ( .D(D_19), .E(n6431), .C(wclk), .QN(n5885) );
  DFE1 \mem_reg_10][18  ( .D(D_18), .E(n6431), .C(wclk), .QN(n5886) );
  DFE1 \mem_reg_10][17  ( .D(D_17), .E(n6431), .C(wclk), .QN(n5887) );
  DFE1 \mem_reg_10][16  ( .D(D_16), .E(n6431), .C(wclk), .QN(n5888) );
  DFE1 \mem_reg_10][15  ( .D(D_15), .E(n6431), .C(wclk), .QN(n5889) );
  DFE1 \mem_reg_10][14  ( .D(D_14), .E(n6431), .C(wclk), .QN(n5890) );
  DFE1 \mem_reg_10][13  ( .D(D_13), .E(n6431), .C(wclk), .QN(n5891) );
  DFE1 \mem_reg_10][12  ( .D(D_12), .E(n6431), .C(wclk), .QN(n5892) );
  DFE1 \mem_reg_10][11  ( .D(D_11), .E(n6431), .C(wclk), .QN(n5893) );
  DFE1 \mem_reg_10][10  ( .D(D_10), .E(n6431), .C(wclk), .QN(n5894) );
  DFE1 \mem_reg_10][9  ( .D(D_9), .E(n6431), .C(wclk), .QN(n5895) );
  DFE1 \mem_reg_10][8  ( .D(D_8), .E(n6431), .C(wclk), .QN(n5896) );
  DFE1 \mem_reg_10][7  ( .D(D_7), .E(n6431), .C(wclk), .QN(n5897) );
  DFE1 \mem_reg_10][6  ( .D(D_6), .E(n6431), .C(wclk), .QN(n5898) );
  DFE1 \mem_reg_10][5  ( .D(D_5), .E(n6431), .C(wclk), .QN(n5899) );
  DFE1 \mem_reg_10][4  ( .D(D_4), .E(n6431), .C(wclk), .QN(n5900) );
  DFE1 \mem_reg_10][3  ( .D(D_3), .E(n6431), .C(wclk), .QN(n5901) );
  DFE1 \mem_reg_10][2  ( .D(D_2), .E(n6431), .C(wclk), .QN(n5902) );
  DFE1 \mem_reg_10][1  ( .D(D_1), .E(n6431), .C(wclk), .QN(n5903) );
  DFE1 \mem_reg_10][0  ( .D(D_0), .E(n6431), .C(wclk), .QN(n5904) );
  DFE1 \mem_reg_55][23  ( .D(D_23), .E(n6490), .C(wclk), .QN(n4801) );
  DFE1 \mem_reg_55][22  ( .D(D_22), .E(n6490), .C(wclk), .QN(n4802) );
  DFE1 \mem_reg_55][21  ( .D(D_21), .E(n6490), .C(wclk), .QN(n4803) );
  DFE1 \mem_reg_55][20  ( .D(D_20), .E(n6490), .C(wclk), .QN(n4804) );
  DFE1 \mem_reg_55][19  ( .D(D_19), .E(n6490), .C(wclk), .QN(n4805) );
  DFE1 \mem_reg_55][18  ( .D(D_18), .E(n6490), .C(wclk), .QN(n4806) );
  DFE1 \mem_reg_55][17  ( .D(D_17), .E(n6490), .C(wclk), .QN(n4807) );
  DFE1 \mem_reg_55][16  ( .D(D_16), .E(n6490), .C(wclk), .QN(n4808) );
  DFE1 \mem_reg_55][15  ( .D(D_15), .E(n6490), .C(wclk), .QN(n4809) );
  DFE1 \mem_reg_55][14  ( .D(D_14), .E(n6490), .C(wclk), .QN(n4810) );
  DFE1 \mem_reg_55][13  ( .D(D_13), .E(n6490), .C(wclk), .QN(n4811) );
  DFE1 \mem_reg_55][12  ( .D(D_12), .E(n6490), .C(wclk), .QN(n4812) );
  DFE1 \mem_reg_55][11  ( .D(D_11), .E(n6490), .C(wclk), .QN(n4813) );
  DFE1 \mem_reg_55][10  ( .D(D_10), .E(n6490), .C(wclk), .QN(n4814) );
  DFE1 \mem_reg_55][9  ( .D(D_9), .E(n6490), .C(wclk), .QN(n4815) );
  DFE1 \mem_reg_55][8  ( .D(D_8), .E(n6490), .C(wclk), .QN(n4816) );
  DFE1 \mem_reg_55][7  ( .D(D_7), .E(n6490), .C(wclk), .QN(n4817) );
  DFE1 \mem_reg_55][6  ( .D(D_6), .E(n6490), .C(wclk), .QN(n4818) );
  DFE1 \mem_reg_55][5  ( .D(D_5), .E(n6490), .C(wclk), .QN(n4819) );
  DFE1 \mem_reg_55][4  ( .D(D_4), .E(n6490), .C(wclk), .QN(n4820) );
  DFE1 \mem_reg_55][3  ( .D(D_3), .E(n6490), .C(wclk), .QN(n4821) );
  DFE1 \mem_reg_55][2  ( .D(D_2), .E(n6490), .C(wclk), .QN(n4822) );
  DFE1 \mem_reg_55][1  ( .D(D_1), .E(n6490), .C(wclk), .QN(n4823) );
  DFE1 \mem_reg_55][0  ( .D(D_0), .E(n6490), .C(wclk), .QN(n4824) );
  DFE1 \mem_reg_54][23  ( .D(D_23), .E(n6489), .C(wclk), .QN(n4825) );
  DFE1 \mem_reg_54][22  ( .D(D_22), .E(n6489), .C(wclk), .QN(n4826) );
  DFE1 \mem_reg_54][21  ( .D(D_21), .E(n6489), .C(wclk), .QN(n4827) );
  DFE1 \mem_reg_54][20  ( .D(D_20), .E(n6489), .C(wclk), .QN(n4828) );
  DFE1 \mem_reg_54][19  ( .D(D_19), .E(n6489), .C(wclk), .QN(n4829) );
  DFE1 \mem_reg_54][18  ( .D(D_18), .E(n6489), .C(wclk), .QN(n4830) );
  DFE1 \mem_reg_54][17  ( .D(D_17), .E(n6489), .C(wclk), .QN(n4831) );
  DFE1 \mem_reg_54][16  ( .D(D_16), .E(n6489), .C(wclk), .QN(n4832) );
  DFE1 \mem_reg_54][15  ( .D(D_15), .E(n6489), .C(wclk), .QN(n4833) );
  DFE1 \mem_reg_54][14  ( .D(D_14), .E(n6489), .C(wclk), .QN(n4834) );
  DFE1 \mem_reg_54][13  ( .D(D_13), .E(n6489), .C(wclk), .QN(n4835) );
  DFE1 \mem_reg_54][12  ( .D(D_12), .E(n6489), .C(wclk), .QN(n4836) );
  DFE1 \mem_reg_54][11  ( .D(D_11), .E(n6489), .C(wclk), .QN(n4837) );
  DFE1 \mem_reg_54][10  ( .D(D_10), .E(n6489), .C(wclk), .QN(n4838) );
  DFE1 \mem_reg_54][9  ( .D(D_9), .E(n6489), .C(wclk), .QN(n4839) );
  DFE1 \mem_reg_54][8  ( .D(D_8), .E(n6489), .C(wclk), .QN(n4840) );
  DFE1 \mem_reg_54][7  ( .D(D_7), .E(n6489), .C(wclk), .QN(n4841) );
  DFE1 \mem_reg_54][6  ( .D(D_6), .E(n6489), .C(wclk), .QN(n4842) );
  DFE1 \mem_reg_54][5  ( .D(D_5), .E(n6489), .C(wclk), .QN(n4843) );
  DFE1 \mem_reg_54][4  ( .D(D_4), .E(n6489), .C(wclk), .QN(n4844) );
  DFE1 \mem_reg_54][3  ( .D(D_3), .E(n6489), .C(wclk), .QN(n4845) );
  DFE1 \mem_reg_54][2  ( .D(D_2), .E(n6489), .C(wclk), .QN(n4846) );
  DFE1 \mem_reg_54][1  ( .D(D_1), .E(n6489), .C(wclk), .QN(n4847) );
  DFE1 \mem_reg_54][0  ( .D(D_0), .E(n6489), .C(wclk), .QN(n4848) );
  DFE1 \mem_reg_51][23  ( .D(D_23), .E(n6485), .C(wclk), .QN(n4897) );
  DFE1 \mem_reg_51][22  ( .D(D_22), .E(n6485), .C(wclk), .QN(n4898) );
  DFE1 \mem_reg_51][21  ( .D(D_21), .E(n6485), .C(wclk), .QN(n4899) );
  DFE1 \mem_reg_51][20  ( .D(D_20), .E(n6485), .C(wclk), .QN(n4900) );
  DFE1 \mem_reg_51][19  ( .D(D_19), .E(n6485), .C(wclk), .QN(n4901) );
  DFE1 \mem_reg_51][18  ( .D(D_18), .E(n6485), .C(wclk), .QN(n4902) );
  DFE1 \mem_reg_51][17  ( .D(D_17), .E(n6485), .C(wclk), .QN(n4903) );
  DFE1 \mem_reg_51][16  ( .D(D_16), .E(n6485), .C(wclk), .QN(n4904) );
  DFE1 \mem_reg_51][15  ( .D(D_15), .E(n6485), .C(wclk), .QN(n4905) );
  DFE1 \mem_reg_51][14  ( .D(D_14), .E(n6485), .C(wclk), .QN(n4906) );
  DFE1 \mem_reg_51][13  ( .D(D_13), .E(n6485), .C(wclk), .QN(n4907) );
  DFE1 \mem_reg_51][12  ( .D(D_12), .E(n6485), .C(wclk), .QN(n4908) );
  DFE1 \mem_reg_51][11  ( .D(D_11), .E(n6485), .C(wclk), .QN(n4909) );
  DFE1 \mem_reg_51][10  ( .D(D_10), .E(n6485), .C(wclk), .QN(n4910) );
  DFE1 \mem_reg_51][9  ( .D(D_9), .E(n6485), .C(wclk), .QN(n4911) );
  DFE1 \mem_reg_51][8  ( .D(D_8), .E(n6485), .C(wclk), .QN(n4912) );
  DFE1 \mem_reg_51][7  ( .D(D_7), .E(n6485), .C(wclk), .QN(n4913) );
  DFE1 \mem_reg_51][6  ( .D(D_6), .E(n6485), .C(wclk), .QN(n4914) );
  DFE1 \mem_reg_51][5  ( .D(D_5), .E(n6485), .C(wclk), .QN(n4915) );
  DFE1 \mem_reg_51][4  ( .D(D_4), .E(n6485), .C(wclk), .QN(n4916) );
  DFE1 \mem_reg_51][3  ( .D(D_3), .E(n6485), .C(wclk), .QN(n4917) );
  DFE1 \mem_reg_51][2  ( .D(D_2), .E(n6485), .C(wclk), .QN(n4918) );
  DFE1 \mem_reg_51][1  ( .D(D_1), .E(n6485), .C(wclk), .QN(n4919) );
  DFE1 \mem_reg_51][0  ( .D(D_0), .E(n6485), .C(wclk), .QN(n4920) );
  DFE1 \mem_reg_50][23  ( .D(D_23), .E(n6484), .C(wclk), .QN(n4921) );
  DFE1 \mem_reg_50][22  ( .D(D_22), .E(n6484), .C(wclk), .QN(n4922) );
  DFE1 \mem_reg_50][21  ( .D(D_21), .E(n6484), .C(wclk), .QN(n4923) );
  DFE1 \mem_reg_50][20  ( .D(D_20), .E(n6484), .C(wclk), .QN(n4924) );
  DFE1 \mem_reg_50][19  ( .D(D_19), .E(n6484), .C(wclk), .QN(n4925) );
  DFE1 \mem_reg_50][18  ( .D(D_18), .E(n6484), .C(wclk), .QN(n4926) );
  DFE1 \mem_reg_50][17  ( .D(D_17), .E(n6484), .C(wclk), .QN(n4927) );
  DFE1 \mem_reg_50][16  ( .D(D_16), .E(n6484), .C(wclk), .QN(n4928) );
  DFE1 \mem_reg_50][15  ( .D(D_15), .E(n6484), .C(wclk), .QN(n4929) );
  DFE1 \mem_reg_50][14  ( .D(D_14), .E(n6484), .C(wclk), .QN(n4930) );
  DFE1 \mem_reg_50][13  ( .D(D_13), .E(n6484), .C(wclk), .QN(n4931) );
  DFE1 \mem_reg_50][12  ( .D(D_12), .E(n6484), .C(wclk), .QN(n4932) );
  DFE1 \mem_reg_50][11  ( .D(D_11), .E(n6484), .C(wclk), .QN(n4933) );
  DFE1 \mem_reg_50][10  ( .D(D_10), .E(n6484), .C(wclk), .QN(n4934) );
  DFE1 \mem_reg_50][9  ( .D(D_9), .E(n6484), .C(wclk), .QN(n4935) );
  DFE1 \mem_reg_50][8  ( .D(D_8), .E(n6484), .C(wclk), .QN(n4936) );
  DFE1 \mem_reg_50][7  ( .D(D_7), .E(n6484), .C(wclk), .QN(n4937) );
  DFE1 \mem_reg_50][6  ( .D(D_6), .E(n6484), .C(wclk), .QN(n4938) );
  DFE1 \mem_reg_50][5  ( .D(D_5), .E(n6484), .C(wclk), .QN(n4939) );
  DFE1 \mem_reg_50][4  ( .D(D_4), .E(n6484), .C(wclk), .QN(n4940) );
  DFE1 \mem_reg_50][3  ( .D(D_3), .E(n6484), .C(wclk), .QN(n4941) );
  DFE1 \mem_reg_50][2  ( .D(D_2), .E(n6484), .C(wclk), .QN(n4942) );
  DFE1 \mem_reg_50][1  ( .D(D_1), .E(n6484), .C(wclk), .QN(n4943) );
  DFE1 \mem_reg_50][0  ( .D(D_0), .E(n6484), .C(wclk), .QN(n4944) );
  DFE1 \mem_reg_63][23  ( .D(D_23), .E(n6198), .C(wclk), .QN(n4609) );
  DFE1 \mem_reg_63][22  ( .D(D_22), .E(n6198), .C(wclk), .QN(n4610) );
  DFE1 \mem_reg_63][21  ( .D(D_21), .E(n6198), .C(wclk), .QN(n4611) );
  DFE1 \mem_reg_63][20  ( .D(D_20), .E(n6198), .C(wclk), .QN(n4612) );
  DFE1 \mem_reg_63][19  ( .D(D_19), .E(n6198), .C(wclk), .QN(n4613) );
  DFE1 \mem_reg_63][18  ( .D(D_18), .E(n6198), .C(wclk), .QN(n4614) );
  DFE1 \mem_reg_63][17  ( .D(D_17), .E(n6198), .C(wclk), .QN(n4615) );
  DFE1 \mem_reg_63][16  ( .D(D_16), .E(n6198), .C(wclk), .QN(n4616) );
  DFE1 \mem_reg_63][15  ( .D(D_15), .E(n6198), .C(wclk), .QN(n4617) );
  DFE1 \mem_reg_63][14  ( .D(D_14), .E(n6198), .C(wclk), .QN(n4618) );
  DFE1 \mem_reg_63][13  ( .D(D_13), .E(n6198), .C(wclk), .QN(n4619) );
  DFE1 \mem_reg_63][12  ( .D(D_12), .E(n6198), .C(wclk), .QN(n4620) );
  DFE1 \mem_reg_63][11  ( .D(D_11), .E(n6198), .C(wclk), .QN(n4621) );
  DFE1 \mem_reg_63][10  ( .D(D_10), .E(n6198), .C(wclk), .QN(n4622) );
  DFE1 \mem_reg_63][9  ( .D(D_9), .E(n6198), .C(wclk), .QN(n4623) );
  DFE1 \mem_reg_63][8  ( .D(D_8), .E(n6198), .C(wclk), .QN(n4624) );
  DFE1 \mem_reg_63][7  ( .D(D_7), .E(n6198), .C(wclk), .QN(n4625) );
  DFE1 \mem_reg_63][6  ( .D(D_6), .E(n6198), .C(wclk), .QN(n4626) );
  DFE1 \mem_reg_63][5  ( .D(D_5), .E(n6198), .C(wclk), .QN(n4627) );
  DFE1 \mem_reg_63][4  ( .D(D_4), .E(n6198), .C(wclk), .QN(n4628) );
  DFE1 \mem_reg_63][3  ( .D(D_3), .E(n6198), .C(wclk), .QN(n4629) );
  DFE1 \mem_reg_63][2  ( .D(D_2), .E(n6198), .C(wclk), .QN(n4630) );
  DFE1 \mem_reg_63][1  ( .D(D_1), .E(n6198), .C(wclk), .QN(n4631) );
  DFE1 \mem_reg_63][0  ( .D(D_0), .E(n6198), .C(wclk), .QN(n4632) );
  DFE1 \mem_reg_62][23  ( .D(D_23), .E(n6195), .C(wclk), .QN(n4633) );
  DFE1 \mem_reg_62][22  ( .D(D_22), .E(n6195), .C(wclk), .QN(n4634) );
  DFE1 \mem_reg_62][21  ( .D(D_21), .E(n6195), .C(wclk), .QN(n4635) );
  DFE1 \mem_reg_62][20  ( .D(D_20), .E(n6195), .C(wclk), .QN(n4636) );
  DFE1 \mem_reg_62][19  ( .D(D_19), .E(n6195), .C(wclk), .QN(n4637) );
  DFE1 \mem_reg_62][18  ( .D(D_18), .E(n6195), .C(wclk), .QN(n4638) );
  DFE1 \mem_reg_62][17  ( .D(D_17), .E(n6195), .C(wclk), .QN(n4639) );
  DFE1 \mem_reg_62][16  ( .D(D_16), .E(n6195), .C(wclk), .QN(n4640) );
  DFE1 \mem_reg_62][15  ( .D(D_15), .E(n6195), .C(wclk), .QN(n4641) );
  DFE1 \mem_reg_62][14  ( .D(D_14), .E(n6195), .C(wclk), .QN(n4642) );
  DFE1 \mem_reg_62][13  ( .D(D_13), .E(n6195), .C(wclk), .QN(n4643) );
  DFE1 \mem_reg_62][12  ( .D(D_12), .E(n6195), .C(wclk), .QN(n4644) );
  DFE1 \mem_reg_62][11  ( .D(D_11), .E(n6195), .C(wclk), .QN(n4645) );
  DFE1 \mem_reg_62][10  ( .D(D_10), .E(n6195), .C(wclk), .QN(n4646) );
  DFE1 \mem_reg_62][9  ( .D(D_9), .E(n6195), .C(wclk), .QN(n4647) );
  DFE1 \mem_reg_62][8  ( .D(D_8), .E(n6195), .C(wclk), .QN(n4648) );
  DFE1 \mem_reg_62][7  ( .D(D_7), .E(n6195), .C(wclk), .QN(n4649) );
  DFE1 \mem_reg_62][6  ( .D(D_6), .E(n6195), .C(wclk), .QN(n4650) );
  DFE1 \mem_reg_62][5  ( .D(D_5), .E(n6195), .C(wclk), .QN(n4651) );
  DFE1 \mem_reg_62][4  ( .D(D_4), .E(n6195), .C(wclk), .QN(n4652) );
  DFE1 \mem_reg_62][3  ( .D(D_3), .E(n6195), .C(wclk), .QN(n4653) );
  DFE1 \mem_reg_62][2  ( .D(D_2), .E(n6195), .C(wclk), .QN(n4654) );
  DFE1 \mem_reg_62][1  ( .D(D_1), .E(n6195), .C(wclk), .QN(n4655) );
  DFE1 \mem_reg_62][0  ( .D(D_0), .E(n6195), .C(wclk), .QN(n4656) );
  DFE1 \mem_reg_60][23  ( .D(D_23), .E(n6496), .C(wclk), .QN(n4681) );
  DFE1 \mem_reg_60][22  ( .D(D_22), .E(n6496), .C(wclk), .QN(n4682) );
  DFE1 \mem_reg_60][21  ( .D(D_21), .E(n6496), .C(wclk), .QN(n4683) );
  DFE1 \mem_reg_60][20  ( .D(D_20), .E(n6496), .C(wclk), .QN(n4684) );
  DFE1 \mem_reg_60][19  ( .D(D_19), .E(n6496), .C(wclk), .QN(n4685) );
  DFE1 \mem_reg_60][18  ( .D(D_18), .E(n6496), .C(wclk), .QN(n4686) );
  DFE1 \mem_reg_60][17  ( .D(D_17), .E(n6496), .C(wclk), .QN(n4687) );
  DFE1 \mem_reg_60][16  ( .D(D_16), .E(n6496), .C(wclk), .QN(n4688) );
  DFE1 \mem_reg_60][15  ( .D(D_15), .E(n6496), .C(wclk), .QN(n4689) );
  DFE1 \mem_reg_60][14  ( .D(D_14), .E(n6496), .C(wclk), .QN(n4690) );
  DFE1 \mem_reg_60][13  ( .D(D_13), .E(n6496), .C(wclk), .QN(n4691) );
  DFE1 \mem_reg_60][12  ( .D(D_12), .E(n6496), .C(wclk), .QN(n4692) );
  DFE1 \mem_reg_60][11  ( .D(D_11), .E(n6496), .C(wclk), .QN(n4693) );
  DFE1 \mem_reg_60][10  ( .D(D_10), .E(n6496), .C(wclk), .QN(n4694) );
  DFE1 \mem_reg_60][9  ( .D(D_9), .E(n6496), .C(wclk), .QN(n4695) );
  DFE1 \mem_reg_60][8  ( .D(D_8), .E(n6496), .C(wclk), .QN(n4696) );
  DFE1 \mem_reg_60][7  ( .D(D_7), .E(n6496), .C(wclk), .QN(n4697) );
  DFE1 \mem_reg_60][6  ( .D(D_6), .E(n6496), .C(wclk), .QN(n4698) );
  DFE1 \mem_reg_60][5  ( .D(D_5), .E(n6496), .C(wclk), .QN(n4699) );
  DFE1 \mem_reg_60][4  ( .D(D_4), .E(n6496), .C(wclk), .QN(n4700) );
  DFE1 \mem_reg_60][3  ( .D(D_3), .E(n6496), .C(wclk), .QN(n4701) );
  DFE1 \mem_reg_60][2  ( .D(D_2), .E(n6496), .C(wclk), .QN(n4702) );
  DFE1 \mem_reg_60][1  ( .D(D_1), .E(n6496), .C(wclk), .QN(n4703) );
  DFE1 \mem_reg_60][0  ( .D(D_0), .E(n6496), .C(wclk), .QN(n4704) );
  DFE1 \mem_reg_56][23  ( .D(D_23), .E(n6491), .C(wclk), .QN(n4777) );
  DFE1 \mem_reg_56][22  ( .D(D_22), .E(n6491), .C(wclk), .QN(n4778) );
  DFE1 \mem_reg_56][21  ( .D(D_21), .E(n6491), .C(wclk), .QN(n4779) );
  DFE1 \mem_reg_56][20  ( .D(D_20), .E(n6491), .C(wclk), .QN(n4780) );
  DFE1 \mem_reg_56][19  ( .D(D_19), .E(n6491), .C(wclk), .QN(n4781) );
  DFE1 \mem_reg_56][18  ( .D(D_18), .E(n6491), .C(wclk), .QN(n4782) );
  DFE1 \mem_reg_56][17  ( .D(D_17), .E(n6491), .C(wclk), .QN(n4783) );
  DFE1 \mem_reg_56][16  ( .D(D_16), .E(n6491), .C(wclk), .QN(n4784) );
  DFE1 \mem_reg_56][15  ( .D(D_15), .E(n6491), .C(wclk), .QN(n4785) );
  DFE1 \mem_reg_56][14  ( .D(D_14), .E(n6491), .C(wclk), .QN(n4786) );
  DFE1 \mem_reg_56][13  ( .D(D_13), .E(n6491), .C(wclk), .QN(n4787) );
  DFE1 \mem_reg_56][12  ( .D(D_12), .E(n6491), .C(wclk), .QN(n4788) );
  DFE1 \mem_reg_56][11  ( .D(D_11), .E(n6491), .C(wclk), .QN(n4789) );
  DFE1 \mem_reg_56][10  ( .D(D_10), .E(n6491), .C(wclk), .QN(n4790) );
  DFE1 \mem_reg_56][9  ( .D(D_9), .E(n6491), .C(wclk), .QN(n4791) );
  DFE1 \mem_reg_56][8  ( .D(D_8), .E(n6491), .C(wclk), .QN(n4792) );
  DFE1 \mem_reg_56][7  ( .D(D_7), .E(n6491), .C(wclk), .QN(n4793) );
  DFE1 \mem_reg_56][6  ( .D(D_6), .E(n6491), .C(wclk), .QN(n4794) );
  DFE1 \mem_reg_56][5  ( .D(D_5), .E(n6491), .C(wclk), .QN(n4795) );
  DFE1 \mem_reg_56][4  ( .D(D_4), .E(n6491), .C(wclk), .QN(n4796) );
  DFE1 \mem_reg_56][3  ( .D(D_3), .E(n6491), .C(wclk), .QN(n4797) );
  DFE1 \mem_reg_56][2  ( .D(D_2), .E(n6491), .C(wclk), .QN(n4798) );
  DFE1 \mem_reg_56][1  ( .D(D_1), .E(n6491), .C(wclk), .QN(n4799) );
  DFE1 \mem_reg_56][0  ( .D(D_0), .E(n6491), .C(wclk), .QN(n4800) );
  DFE1 \mem_reg_52][23  ( .D(D_23), .E(n6486), .C(wclk), .QN(n4873) );
  DFE1 \mem_reg_52][22  ( .D(D_22), .E(n6486), .C(wclk), .QN(n4874) );
  DFE1 \mem_reg_52][21  ( .D(D_21), .E(n6486), .C(wclk), .QN(n4875) );
  DFE1 \mem_reg_52][20  ( .D(D_20), .E(n6486), .C(wclk), .QN(n4876) );
  DFE1 \mem_reg_52][19  ( .D(D_19), .E(n6486), .C(wclk), .QN(n4877) );
  DFE1 \mem_reg_52][18  ( .D(D_18), .E(n6486), .C(wclk), .QN(n4878) );
  DFE1 \mem_reg_52][17  ( .D(D_17), .E(n6486), .C(wclk), .QN(n4879) );
  DFE1 \mem_reg_52][16  ( .D(D_16), .E(n6486), .C(wclk), .QN(n4880) );
  DFE1 \mem_reg_52][15  ( .D(D_15), .E(n6486), .C(wclk), .QN(n4881) );
  DFE1 \mem_reg_52][14  ( .D(D_14), .E(n6486), .C(wclk), .QN(n4882) );
  DFE1 \mem_reg_52][13  ( .D(D_13), .E(n6486), .C(wclk), .QN(n4883) );
  DFE1 \mem_reg_52][12  ( .D(D_12), .E(n6486), .C(wclk), .QN(n4884) );
  DFE1 \mem_reg_52][11  ( .D(D_11), .E(n6486), .C(wclk), .QN(n4885) );
  DFE1 \mem_reg_52][10  ( .D(D_10), .E(n6486), .C(wclk), .QN(n4886) );
  DFE1 \mem_reg_52][9  ( .D(D_9), .E(n6486), .C(wclk), .QN(n4887) );
  DFE1 \mem_reg_52][8  ( .D(D_8), .E(n6486), .C(wclk), .QN(n4888) );
  DFE1 \mem_reg_52][7  ( .D(D_7), .E(n6486), .C(wclk), .QN(n4889) );
  DFE1 \mem_reg_52][6  ( .D(D_6), .E(n6486), .C(wclk), .QN(n4890) );
  DFE1 \mem_reg_52][5  ( .D(D_5), .E(n6486), .C(wclk), .QN(n4891) );
  DFE1 \mem_reg_52][4  ( .D(D_4), .E(n6486), .C(wclk), .QN(n4892) );
  DFE1 \mem_reg_52][3  ( .D(D_3), .E(n6486), .C(wclk), .QN(n4893) );
  DFE1 \mem_reg_52][2  ( .D(D_2), .E(n6486), .C(wclk), .QN(n4894) );
  DFE1 \mem_reg_52][1  ( .D(D_1), .E(n6486), .C(wclk), .QN(n4895) );
  DFE1 \mem_reg_52][0  ( .D(D_0), .E(n6486), .C(wclk), .QN(n4896) );
  DFE1 \mem_reg_48][23  ( .D(D_23), .E(n6479), .C(wclk), .QN(n4969) );
  DFE1 \mem_reg_48][22  ( .D(D_22), .E(n6479), .C(wclk), .QN(n4970) );
  DFE1 \mem_reg_48][21  ( .D(D_21), .E(n6479), .C(wclk), .QN(n4971) );
  DFE1 \mem_reg_48][20  ( .D(D_20), .E(n6479), .C(wclk), .QN(n4972) );
  DFE1 \mem_reg_48][19  ( .D(D_19), .E(n6479), .C(wclk), .QN(n4973) );
  DFE1 \mem_reg_48][18  ( .D(D_18), .E(n6479), .C(wclk), .QN(n4974) );
  DFE1 \mem_reg_48][17  ( .D(D_17), .E(n6479), .C(wclk), .QN(n4975) );
  DFE1 \mem_reg_48][16  ( .D(D_16), .E(n6479), .C(wclk), .QN(n4976) );
  DFE1 \mem_reg_48][15  ( .D(D_15), .E(n6479), .C(wclk), .QN(n4977) );
  DFE1 \mem_reg_48][14  ( .D(D_14), .E(n6479), .C(wclk), .QN(n4978) );
  DFE1 \mem_reg_48][13  ( .D(D_13), .E(n6479), .C(wclk), .QN(n4979) );
  DFE1 \mem_reg_48][12  ( .D(D_12), .E(n6479), .C(wclk), .QN(n4980) );
  DFE1 \mem_reg_48][11  ( .D(D_11), .E(n6479), .C(wclk), .QN(n4981) );
  DFE1 \mem_reg_48][10  ( .D(D_10), .E(n6479), .C(wclk), .QN(n4982) );
  DFE1 \mem_reg_48][9  ( .D(D_9), .E(n6479), .C(wclk), .QN(n4983) );
  DFE1 \mem_reg_48][8  ( .D(D_8), .E(n6479), .C(wclk), .QN(n4984) );
  DFE1 \mem_reg_48][7  ( .D(D_7), .E(n6479), .C(wclk), .QN(n4985) );
  DFE1 \mem_reg_48][6  ( .D(D_6), .E(n6479), .C(wclk), .QN(n4986) );
  DFE1 \mem_reg_48][5  ( .D(D_5), .E(n6479), .C(wclk), .QN(n4987) );
  DFE1 \mem_reg_48][4  ( .D(D_4), .E(n6479), .C(wclk), .QN(n4988) );
  DFE1 \mem_reg_48][3  ( .D(D_3), .E(n6479), .C(wclk), .QN(n4989) );
  DFE1 \mem_reg_48][2  ( .D(D_2), .E(n6479), .C(wclk), .QN(n4990) );
  DFE1 \mem_reg_48][1  ( .D(D_1), .E(n6479), .C(wclk), .QN(n4991) );
  DFE1 \mem_reg_48][0  ( .D(D_0), .E(n6479), .C(wclk), .QN(n4992) );
  DFE1 \mem_reg_57][23  ( .D(D_23), .E(n6492), .C(wclk), .QN(n4753) );
  DFE1 \mem_reg_57][22  ( .D(D_22), .E(n6492), .C(wclk), .QN(n4754) );
  DFE1 \mem_reg_57][21  ( .D(D_21), .E(n6492), .C(wclk), .QN(n4755) );
  DFE1 \mem_reg_57][20  ( .D(D_20), .E(n6492), .C(wclk), .QN(n4756) );
  DFE1 \mem_reg_57][19  ( .D(D_19), .E(n6492), .C(wclk), .QN(n4757) );
  DFE1 \mem_reg_57][18  ( .D(D_18), .E(n6492), .C(wclk), .QN(n4758) );
  DFE1 \mem_reg_57][17  ( .D(D_17), .E(n6492), .C(wclk), .QN(n4759) );
  DFE1 \mem_reg_57][16  ( .D(D_16), .E(n6492), .C(wclk), .QN(n4760) );
  DFE1 \mem_reg_57][15  ( .D(D_15), .E(n6492), .C(wclk), .QN(n4761) );
  DFE1 \mem_reg_57][14  ( .D(D_14), .E(n6492), .C(wclk), .QN(n4762) );
  DFE1 \mem_reg_57][13  ( .D(D_13), .E(n6492), .C(wclk), .QN(n4763) );
  DFE1 \mem_reg_57][12  ( .D(D_12), .E(n6492), .C(wclk), .QN(n4764) );
  DFE1 \mem_reg_57][11  ( .D(D_11), .E(n6492), .C(wclk), .QN(n4765) );
  DFE1 \mem_reg_57][10  ( .D(D_10), .E(n6492), .C(wclk), .QN(n4766) );
  DFE1 \mem_reg_57][9  ( .D(D_9), .E(n6492), .C(wclk), .QN(n4767) );
  DFE1 \mem_reg_57][8  ( .D(D_8), .E(n6492), .C(wclk), .QN(n4768) );
  DFE1 \mem_reg_57][7  ( .D(D_7), .E(n6492), .C(wclk), .QN(n4769) );
  DFE1 \mem_reg_57][6  ( .D(D_6), .E(n6492), .C(wclk), .QN(n4770) );
  DFE1 \mem_reg_57][5  ( .D(D_5), .E(n6492), .C(wclk), .QN(n4771) );
  DFE1 \mem_reg_57][4  ( .D(D_4), .E(n6492), .C(wclk), .QN(n4772) );
  DFE1 \mem_reg_57][3  ( .D(D_3), .E(n6492), .C(wclk), .QN(n4773) );
  DFE1 \mem_reg_57][2  ( .D(D_2), .E(n6492), .C(wclk), .QN(n4774) );
  DFE1 \mem_reg_57][1  ( .D(D_1), .E(n6492), .C(wclk), .QN(n4775) );
  DFE1 \mem_reg_57][0  ( .D(D_0), .E(n6492), .C(wclk), .QN(n4776) );
  DFE1 \mem_reg_53][23  ( .D(D_23), .E(n6488), .C(wclk), .QN(n4849) );
  DFE1 \mem_reg_53][22  ( .D(D_22), .E(n6488), .C(wclk), .QN(n4850) );
  DFE1 \mem_reg_53][21  ( .D(D_21), .E(n6488), .C(wclk), .QN(n4851) );
  DFE1 \mem_reg_53][20  ( .D(D_20), .E(n6488), .C(wclk), .QN(n4852) );
  DFE1 \mem_reg_53][19  ( .D(D_19), .E(n6488), .C(wclk), .QN(n4853) );
  DFE1 \mem_reg_53][18  ( .D(D_18), .E(n6488), .C(wclk), .QN(n4854) );
  DFE1 \mem_reg_53][17  ( .D(D_17), .E(n6488), .C(wclk), .QN(n4855) );
  DFE1 \mem_reg_53][16  ( .D(D_16), .E(n6488), .C(wclk), .QN(n4856) );
  DFE1 \mem_reg_53][15  ( .D(D_15), .E(n6488), .C(wclk), .QN(n4857) );
  DFE1 \mem_reg_53][14  ( .D(D_14), .E(n6488), .C(wclk), .QN(n4858) );
  DFE1 \mem_reg_53][13  ( .D(D_13), .E(n6488), .C(wclk), .QN(n4859) );
  DFE1 \mem_reg_53][12  ( .D(D_12), .E(n6488), .C(wclk), .QN(n4860) );
  DFE1 \mem_reg_53][11  ( .D(D_11), .E(n6488), .C(wclk), .QN(n4861) );
  DFE1 \mem_reg_53][10  ( .D(D_10), .E(n6488), .C(wclk), .QN(n4862) );
  DFE1 \mem_reg_53][9  ( .D(D_9), .E(n6488), .C(wclk), .QN(n4863) );
  DFE1 \mem_reg_53][8  ( .D(D_8), .E(n6488), .C(wclk), .QN(n4864) );
  DFE1 \mem_reg_53][7  ( .D(D_7), .E(n6488), .C(wclk), .QN(n4865) );
  DFE1 \mem_reg_53][6  ( .D(D_6), .E(n6488), .C(wclk), .QN(n4866) );
  DFE1 \mem_reg_53][5  ( .D(D_5), .E(n6488), .C(wclk), .QN(n4867) );
  DFE1 \mem_reg_53][4  ( .D(D_4), .E(n6488), .C(wclk), .QN(n4868) );
  DFE1 \mem_reg_53][3  ( .D(D_3), .E(n6488), .C(wclk), .QN(n4869) );
  DFE1 \mem_reg_53][2  ( .D(D_2), .E(n6488), .C(wclk), .QN(n4870) );
  DFE1 \mem_reg_53][1  ( .D(D_1), .E(n6488), .C(wclk), .QN(n4871) );
  DFE1 \mem_reg_53][0  ( .D(D_0), .E(n6488), .C(wclk), .QN(n4872) );
  DFE1 \mem_reg_49][23  ( .D(D_23), .E(n6482), .C(wclk), .QN(n4945) );
  DFE1 \mem_reg_49][22  ( .D(D_22), .E(n6482), .C(wclk), .QN(n4946) );
  DFE1 \mem_reg_49][21  ( .D(D_21), .E(n6482), .C(wclk), .QN(n4947) );
  DFE1 \mem_reg_49][20  ( .D(D_20), .E(n6482), .C(wclk), .QN(n4948) );
  DFE1 \mem_reg_49][19  ( .D(D_19), .E(n6482), .C(wclk), .QN(n4949) );
  DFE1 \mem_reg_49][18  ( .D(D_18), .E(n6482), .C(wclk), .QN(n4950) );
  DFE1 \mem_reg_49][17  ( .D(D_17), .E(n6482), .C(wclk), .QN(n4951) );
  DFE1 \mem_reg_49][16  ( .D(D_16), .E(n6482), .C(wclk), .QN(n4952) );
  DFE1 \mem_reg_49][15  ( .D(D_15), .E(n6482), .C(wclk), .QN(n4953) );
  DFE1 \mem_reg_49][14  ( .D(D_14), .E(n6482), .C(wclk), .QN(n4954) );
  DFE1 \mem_reg_49][13  ( .D(D_13), .E(n6482), .C(wclk), .QN(n4955) );
  DFE1 \mem_reg_49][12  ( .D(D_12), .E(n6482), .C(wclk), .QN(n4956) );
  DFE1 \mem_reg_49][11  ( .D(D_11), .E(n6482), .C(wclk), .QN(n4957) );
  DFE1 \mem_reg_49][10  ( .D(D_10), .E(n6482), .C(wclk), .QN(n4958) );
  DFE1 \mem_reg_49][9  ( .D(D_9), .E(n6482), .C(wclk), .QN(n4959) );
  DFE1 \mem_reg_49][8  ( .D(D_8), .E(n6482), .C(wclk), .QN(n4960) );
  DFE1 \mem_reg_49][7  ( .D(D_7), .E(n6482), .C(wclk), .QN(n4961) );
  DFE1 \mem_reg_49][6  ( .D(D_6), .E(n6482), .C(wclk), .QN(n4962) );
  DFE1 \mem_reg_49][5  ( .D(D_5), .E(n6482), .C(wclk), .QN(n4963) );
  DFE1 \mem_reg_49][4  ( .D(D_4), .E(n6482), .C(wclk), .QN(n4964) );
  DFE1 \mem_reg_49][3  ( .D(D_3), .E(n6482), .C(wclk), .QN(n4965) );
  DFE1 \mem_reg_49][2  ( .D(D_2), .E(n6482), .C(wclk), .QN(n4966) );
  DFE1 \mem_reg_49][1  ( .D(D_1), .E(n6482), .C(wclk), .QN(n4967) );
  DFE1 \mem_reg_49][0  ( .D(D_0), .E(n6482), .C(wclk), .QN(n4968) );
  DFE1 \mem_reg_13][23  ( .D(D_23), .E(n6434), .C(wclk), .QN(n5809) );
  DFE1 \mem_reg_13][22  ( .D(D_22), .E(n6434), .C(wclk), .QN(n5810) );
  DFE1 \mem_reg_13][21  ( .D(D_21), .E(n6434), .C(wclk), .QN(n5811) );
  DFE1 \mem_reg_13][20  ( .D(D_20), .E(n6434), .C(wclk), .QN(n5812) );
  DFE1 \mem_reg_13][19  ( .D(D_19), .E(n6434), .C(wclk), .QN(n5813) );
  DFE1 \mem_reg_13][18  ( .D(D_18), .E(n6434), .C(wclk), .QN(n5814) );
  DFE1 \mem_reg_13][17  ( .D(D_17), .E(n6434), .C(wclk), .QN(n5815) );
  DFE1 \mem_reg_13][16  ( .D(D_16), .E(n6434), .C(wclk), .QN(n5816) );
  DFE1 \mem_reg_13][15  ( .D(D_15), .E(n6434), .C(wclk), .QN(n5817) );
  DFE1 \mem_reg_13][14  ( .D(D_14), .E(n6434), .C(wclk), .QN(n5818) );
  DFE1 \mem_reg_13][13  ( .D(D_13), .E(n6434), .C(wclk), .QN(n5819) );
  DFE1 \mem_reg_13][12  ( .D(D_12), .E(n6434), .C(wclk), .QN(n5820) );
  DFE1 \mem_reg_13][11  ( .D(D_11), .E(n6434), .C(wclk), .QN(n5821) );
  DFE1 \mem_reg_13][10  ( .D(D_10), .E(n6434), .C(wclk), .QN(n5822) );
  DFE1 \mem_reg_13][9  ( .D(D_9), .E(n6434), .C(wclk), .QN(n5823) );
  DFE1 \mem_reg_13][8  ( .D(D_8), .E(n6434), .C(wclk), .QN(n5824) );
  DFE1 \mem_reg_13][7  ( .D(D_7), .E(n6434), .C(wclk), .QN(n5825) );
  DFE1 \mem_reg_13][6  ( .D(D_6), .E(n6434), .C(wclk), .QN(n5826) );
  DFE1 \mem_reg_13][5  ( .D(D_5), .E(n6434), .C(wclk), .QN(n5827) );
  DFE1 \mem_reg_13][4  ( .D(D_4), .E(n6434), .C(wclk), .QN(n5828) );
  DFE1 \mem_reg_13][3  ( .D(D_3), .E(n6434), .C(wclk), .QN(n5829) );
  DFE1 \mem_reg_13][2  ( .D(D_2), .E(n6434), .C(wclk), .QN(n5830) );
  DFE1 \mem_reg_13][1  ( .D(D_1), .E(n6434), .C(wclk), .QN(n5831) );
  DFE1 \mem_reg_13][0  ( .D(D_0), .E(n6434), .C(wclk), .QN(n5832) );
  DFE1 \mem_reg_5][23  ( .D(D_23), .E(n6426), .C(wclk), .QN(n6001) );
  DFE1 \mem_reg_5][22  ( .D(D_22), .E(n6426), .C(wclk), .QN(n6002) );
  DFE1 \mem_reg_5][21  ( .D(D_21), .E(n6426), .C(wclk), .QN(n6003) );
  DFE1 \mem_reg_5][20  ( .D(D_20), .E(n6426), .C(wclk), .QN(n6004) );
  DFE1 \mem_reg_5][19  ( .D(D_19), .E(n6426), .C(wclk), .QN(n6005) );
  DFE1 \mem_reg_5][18  ( .D(D_18), .E(n6426), .C(wclk), .QN(n6006) );
  DFE1 \mem_reg_5][17  ( .D(D_17), .E(n6426), .C(wclk), .QN(n6007) );
  DFE1 \mem_reg_5][16  ( .D(D_16), .E(n6426), .C(wclk), .QN(n6008) );
  DFE1 \mem_reg_5][15  ( .D(D_15), .E(n6426), .C(wclk), .QN(n6009) );
  DFE1 \mem_reg_5][14  ( .D(D_14), .E(n6426), .C(wclk), .QN(n6010) );
  DFE1 \mem_reg_5][13  ( .D(D_13), .E(n6426), .C(wclk), .QN(n6011) );
  DFE1 \mem_reg_5][12  ( .D(D_12), .E(n6426), .C(wclk), .QN(n6012) );
  DFE1 \mem_reg_5][11  ( .D(D_11), .E(n6426), .C(wclk), .QN(n6013) );
  DFE1 \mem_reg_5][10  ( .D(D_10), .E(n6426), .C(wclk), .QN(n6014) );
  DFE1 \mem_reg_5][9  ( .D(D_9), .E(n6426), .C(wclk), .QN(n6015) );
  DFE1 \mem_reg_5][8  ( .D(D_8), .E(n6426), .C(wclk), .QN(n6016) );
  DFE1 \mem_reg_5][7  ( .D(D_7), .E(n6426), .C(wclk), .QN(n6017) );
  DFE1 \mem_reg_5][6  ( .D(D_6), .E(n6426), .C(wclk), .QN(n6018) );
  DFE1 \mem_reg_5][5  ( .D(D_5), .E(n6426), .C(wclk), .QN(n6019) );
  DFE1 \mem_reg_5][4  ( .D(D_4), .E(n6426), .C(wclk), .QN(n6020) );
  DFE1 \mem_reg_5][3  ( .D(D_3), .E(n6426), .C(wclk), .QN(n6021) );
  DFE1 \mem_reg_5][2  ( .D(D_2), .E(n6426), .C(wclk), .QN(n6022) );
  DFE1 \mem_reg_5][1  ( .D(D_1), .E(n6426), .C(wclk), .QN(n6023) );
  DFE1 \mem_reg_5][0  ( .D(D_0), .E(n6426), .C(wclk), .QN(n6024) );
  DFE1 \mem_reg_1][23  ( .D(D_23), .E(n6421), .C(wclk), .QN(n6097) );
  DFE1 \mem_reg_1][22  ( .D(D_22), .E(n6421), .C(wclk), .QN(n6098) );
  DFE1 \mem_reg_1][21  ( .D(D_21), .E(n6421), .C(wclk), .QN(n6099) );
  DFE1 \mem_reg_1][20  ( .D(D_20), .E(n6421), .C(wclk), .QN(n6100) );
  DFE1 \mem_reg_1][19  ( .D(D_19), .E(n6421), .C(wclk), .QN(n6101) );
  DFE1 \mem_reg_1][18  ( .D(D_18), .E(n6421), .C(wclk), .QN(n6102) );
  DFE1 \mem_reg_1][17  ( .D(D_17), .E(n6421), .C(wclk), .QN(n6103) );
  DFE1 \mem_reg_1][16  ( .D(D_16), .E(n6421), .C(wclk), .QN(n6104) );
  DFE1 \mem_reg_1][15  ( .D(D_15), .E(n6421), .C(wclk), .QN(n6105) );
  DFE1 \mem_reg_1][14  ( .D(D_14), .E(n6421), .C(wclk), .QN(n6106) );
  DFE1 \mem_reg_1][13  ( .D(D_13), .E(n6421), .C(wclk), .QN(n6107) );
  DFE1 \mem_reg_1][12  ( .D(D_12), .E(n6421), .C(wclk), .QN(n6108) );
  DFE1 \mem_reg_1][11  ( .D(D_11), .E(n6421), .C(wclk), .QN(n6109) );
  DFE1 \mem_reg_1][10  ( .D(D_10), .E(n6421), .C(wclk), .QN(n6110) );
  DFE1 \mem_reg_1][9  ( .D(D_9), .E(n6421), .C(wclk), .QN(n6111) );
  DFE1 \mem_reg_1][8  ( .D(D_8), .E(n6421), .C(wclk), .QN(n6112) );
  DFE1 \mem_reg_1][7  ( .D(D_7), .E(n6421), .C(wclk), .QN(n6113) );
  DFE1 \mem_reg_1][6  ( .D(D_6), .E(n6421), .C(wclk), .QN(n6114) );
  DFE1 \mem_reg_1][5  ( .D(D_5), .E(n6421), .C(wclk), .QN(n6115) );
  DFE1 \mem_reg_1][4  ( .D(D_4), .E(n6421), .C(wclk), .QN(n6116) );
  DFE1 \mem_reg_1][3  ( .D(D_3), .E(n6421), .C(wclk), .QN(n6117) );
  DFE1 \mem_reg_1][2  ( .D(D_2), .E(n6421), .C(wclk), .QN(n6118) );
  DFE1 \mem_reg_1][1  ( .D(D_1), .E(n6421), .C(wclk), .QN(n6119) );
  DFE1 \mem_reg_1][0  ( .D(D_0), .E(n6421), .C(wclk), .QN(n6120) );
  DFE1 \mem_reg_207][23  ( .D(D_23), .E(n6380), .C(wclk), .QN(n1153) );
  DFE1 \mem_reg_207][22  ( .D(D_22), .E(n6380), .C(wclk), .QN(n1154) );
  DFE1 \mem_reg_207][21  ( .D(D_21), .E(n6380), .C(wclk), .QN(n1155) );
  DFE1 \mem_reg_207][20  ( .D(D_20), .E(n6380), .C(wclk), .QN(n1156) );
  DFE1 \mem_reg_207][19  ( .D(D_19), .E(n6380), .C(wclk), .QN(n1157) );
  DFE1 \mem_reg_207][18  ( .D(D_18), .E(n6380), .C(wclk), .QN(n1158) );
  DFE1 \mem_reg_207][17  ( .D(D_17), .E(n6380), .C(wclk), .QN(n1159) );
  DFE1 \mem_reg_207][16  ( .D(D_16), .E(n6380), .C(wclk), .QN(n1160) );
  DFE1 \mem_reg_207][15  ( .D(D_15), .E(n6380), .C(wclk), .QN(n1161) );
  DFE1 \mem_reg_207][14  ( .D(D_14), .E(n6380), .C(wclk), .QN(n1162) );
  DFE1 \mem_reg_207][13  ( .D(D_13), .E(n6380), .C(wclk), .QN(n1163) );
  DFE1 \mem_reg_207][12  ( .D(D_12), .E(n6380), .C(wclk), .QN(n1164) );
  DFE1 \mem_reg_207][11  ( .D(D_11), .E(n6380), .C(wclk), .QN(n1165) );
  DFE1 \mem_reg_207][10  ( .D(D_10), .E(n6380), .C(wclk), .QN(n1166) );
  DFE1 \mem_reg_207][9  ( .D(D_9), .E(n6380), .C(wclk), .QN(n1167) );
  DFE1 \mem_reg_207][8  ( .D(D_8), .E(n6380), .C(wclk), .QN(n1168) );
  DFE1 \mem_reg_207][7  ( .D(D_7), .E(n6380), .C(wclk), .QN(n1169) );
  DFE1 \mem_reg_207][6  ( .D(D_6), .E(n6380), .C(wclk), .QN(n1170) );
  DFE1 \mem_reg_207][5  ( .D(D_5), .E(n6380), .C(wclk), .QN(n1171) );
  DFE1 \mem_reg_207][4  ( .D(D_4), .E(n6380), .C(wclk), .QN(n1172) );
  DFE1 \mem_reg_207][3  ( .D(D_3), .E(n6380), .C(wclk), .QN(n1173) );
  DFE1 \mem_reg_207][2  ( .D(D_2), .E(n6380), .C(wclk), .QN(n1174) );
  DFE1 \mem_reg_207][1  ( .D(D_1), .E(n6380), .C(wclk), .QN(n1175) );
  DFE1 \mem_reg_207][0  ( .D(D_0), .E(n6380), .C(wclk), .QN(n1176) );
  DFE1 \mem_reg_206][23  ( .D(D_23), .E(n6379), .C(wclk), .QN(n1177) );
  DFE1 \mem_reg_206][22  ( .D(D_22), .E(n6379), .C(wclk), .QN(n1178) );
  DFE1 \mem_reg_206][21  ( .D(D_21), .E(n6379), .C(wclk), .QN(n1179) );
  DFE1 \mem_reg_206][20  ( .D(D_20), .E(n6379), .C(wclk), .QN(n1180) );
  DFE1 \mem_reg_206][19  ( .D(D_19), .E(n6379), .C(wclk), .QN(n1181) );
  DFE1 \mem_reg_206][18  ( .D(D_18), .E(n6379), .C(wclk), .QN(n1182) );
  DFE1 \mem_reg_206][17  ( .D(D_17), .E(n6379), .C(wclk), .QN(n1183) );
  DFE1 \mem_reg_206][16  ( .D(D_16), .E(n6379), .C(wclk), .QN(n1184) );
  DFE1 \mem_reg_206][15  ( .D(D_15), .E(n6379), .C(wclk), .QN(n1185) );
  DFE1 \mem_reg_206][14  ( .D(D_14), .E(n6379), .C(wclk), .QN(n1186) );
  DFE1 \mem_reg_206][13  ( .D(D_13), .E(n6379), .C(wclk), .QN(n1187) );
  DFE1 \mem_reg_206][12  ( .D(D_12), .E(n6379), .C(wclk), .QN(n1188) );
  DFE1 \mem_reg_206][11  ( .D(D_11), .E(n6379), .C(wclk), .QN(n1189) );
  DFE1 \mem_reg_206][10  ( .D(D_10), .E(n6379), .C(wclk), .QN(n1190) );
  DFE1 \mem_reg_206][9  ( .D(D_9), .E(n6379), .C(wclk), .QN(n1191) );
  DFE1 \mem_reg_206][8  ( .D(D_8), .E(n6379), .C(wclk), .QN(n1192) );
  DFE1 \mem_reg_206][7  ( .D(D_7), .E(n6379), .C(wclk), .QN(n1193) );
  DFE1 \mem_reg_206][6  ( .D(D_6), .E(n6379), .C(wclk), .QN(n1194) );
  DFE1 \mem_reg_206][5  ( .D(D_5), .E(n6379), .C(wclk), .QN(n1195) );
  DFE1 \mem_reg_206][4  ( .D(D_4), .E(n6379), .C(wclk), .QN(n1196) );
  DFE1 \mem_reg_206][3  ( .D(D_3), .E(n6379), .C(wclk), .QN(n1197) );
  DFE1 \mem_reg_206][2  ( .D(D_2), .E(n6379), .C(wclk), .QN(n1198) );
  DFE1 \mem_reg_206][1  ( .D(D_1), .E(n6379), .C(wclk), .QN(n1199) );
  DFE1 \mem_reg_206][0  ( .D(D_0), .E(n6379), .C(wclk), .QN(n1200) );
  DFE1 \mem_reg_205][23  ( .D(D_23), .E(n6378), .C(wclk), .QN(n1201) );
  DFE1 \mem_reg_205][22  ( .D(D_22), .E(n6378), .C(wclk), .QN(n1202) );
  DFE1 \mem_reg_205][21  ( .D(D_21), .E(n6378), .C(wclk), .QN(n1203) );
  DFE1 \mem_reg_205][20  ( .D(D_20), .E(n6378), .C(wclk), .QN(n1204) );
  DFE1 \mem_reg_205][19  ( .D(D_19), .E(n6378), .C(wclk), .QN(n1205) );
  DFE1 \mem_reg_205][18  ( .D(D_18), .E(n6378), .C(wclk), .QN(n1206) );
  DFE1 \mem_reg_205][17  ( .D(D_17), .E(n6378), .C(wclk), .QN(n1207) );
  DFE1 \mem_reg_205][16  ( .D(D_16), .E(n6378), .C(wclk), .QN(n1208) );
  DFE1 \mem_reg_205][15  ( .D(D_15), .E(n6378), .C(wclk), .QN(n1209) );
  DFE1 \mem_reg_205][14  ( .D(D_14), .E(n6378), .C(wclk), .QN(n1210) );
  DFE1 \mem_reg_205][13  ( .D(D_13), .E(n6378), .C(wclk), .QN(n1211) );
  DFE1 \mem_reg_205][12  ( .D(D_12), .E(n6378), .C(wclk), .QN(n1212) );
  DFE1 \mem_reg_205][11  ( .D(D_11), .E(n6378), .C(wclk), .QN(n1213) );
  DFE1 \mem_reg_205][10  ( .D(D_10), .E(n6378), .C(wclk), .QN(n1214) );
  DFE1 \mem_reg_205][9  ( .D(D_9), .E(n6378), .C(wclk), .QN(n1215) );
  DFE1 \mem_reg_205][8  ( .D(D_8), .E(n6378), .C(wclk), .QN(n1216) );
  DFE1 \mem_reg_205][7  ( .D(D_7), .E(n6378), .C(wclk), .QN(n1217) );
  DFE1 \mem_reg_205][6  ( .D(D_6), .E(n6378), .C(wclk), .QN(n1218) );
  DFE1 \mem_reg_205][5  ( .D(D_5), .E(n6378), .C(wclk), .QN(n1219) );
  DFE1 \mem_reg_205][4  ( .D(D_4), .E(n6378), .C(wclk), .QN(n1220) );
  DFE1 \mem_reg_205][3  ( .D(D_3), .E(n6378), .C(wclk), .QN(n1221) );
  DFE1 \mem_reg_205][2  ( .D(D_2), .E(n6378), .C(wclk), .QN(n1222) );
  DFE1 \mem_reg_205][1  ( .D(D_1), .E(n6378), .C(wclk), .QN(n1223) );
  DFE1 \mem_reg_205][0  ( .D(D_0), .E(n6378), .C(wclk), .QN(n1224) );
  DFE1 \mem_reg_204][23  ( .D(D_23), .E(n6377), .C(wclk), .QN(n1225) );
  DFE1 \mem_reg_204][22  ( .D(D_22), .E(n6377), .C(wclk), .QN(n1226) );
  DFE1 \mem_reg_204][21  ( .D(D_21), .E(n6377), .C(wclk), .QN(n1227) );
  DFE1 \mem_reg_204][20  ( .D(D_20), .E(n6377), .C(wclk), .QN(n1228) );
  DFE1 \mem_reg_204][19  ( .D(D_19), .E(n6377), .C(wclk), .QN(n1229) );
  DFE1 \mem_reg_204][18  ( .D(D_18), .E(n6377), .C(wclk), .QN(n1230) );
  DFE1 \mem_reg_204][17  ( .D(D_17), .E(n6377), .C(wclk), .QN(n1231) );
  DFE1 \mem_reg_204][16  ( .D(D_16), .E(n6377), .C(wclk), .QN(n1232) );
  DFE1 \mem_reg_204][15  ( .D(D_15), .E(n6377), .C(wclk), .QN(n1233) );
  DFE1 \mem_reg_204][14  ( .D(D_14), .E(n6377), .C(wclk), .QN(n1234) );
  DFE1 \mem_reg_204][13  ( .D(D_13), .E(n6377), .C(wclk), .QN(n1235) );
  DFE1 \mem_reg_204][12  ( .D(D_12), .E(n6377), .C(wclk), .QN(n1236) );
  DFE1 \mem_reg_204][11  ( .D(D_11), .E(n6377), .C(wclk), .QN(n1237) );
  DFE1 \mem_reg_204][10  ( .D(D_10), .E(n6377), .C(wclk), .QN(n1238) );
  DFE1 \mem_reg_204][9  ( .D(D_9), .E(n6377), .C(wclk), .QN(n1239) );
  DFE1 \mem_reg_204][8  ( .D(D_8), .E(n6377), .C(wclk), .QN(n1240) );
  DFE1 \mem_reg_204][7  ( .D(D_7), .E(n6377), .C(wclk), .QN(n1241) );
  DFE1 \mem_reg_204][6  ( .D(D_6), .E(n6377), .C(wclk), .QN(n1242) );
  DFE1 \mem_reg_204][5  ( .D(D_5), .E(n6377), .C(wclk), .QN(n1243) );
  DFE1 \mem_reg_204][4  ( .D(D_4), .E(n6377), .C(wclk), .QN(n1244) );
  DFE1 \mem_reg_204][3  ( .D(D_3), .E(n6377), .C(wclk), .QN(n1245) );
  DFE1 \mem_reg_204][2  ( .D(D_2), .E(n6377), .C(wclk), .QN(n1246) );
  DFE1 \mem_reg_204][1  ( .D(D_1), .E(n6377), .C(wclk), .QN(n1247) );
  DFE1 \mem_reg_204][0  ( .D(D_0), .E(n6377), .C(wclk), .QN(n1248) );
  DFE1 \mem_reg_203][23  ( .D(D_23), .E(n6376), .C(wclk), .QN(n1249) );
  DFE1 \mem_reg_203][22  ( .D(D_22), .E(n6376), .C(wclk), .QN(n1250) );
  DFE1 \mem_reg_203][21  ( .D(D_21), .E(n6376), .C(wclk), .QN(n1251) );
  DFE1 \mem_reg_203][20  ( .D(D_20), .E(n6376), .C(wclk), .QN(n1252) );
  DFE1 \mem_reg_203][19  ( .D(D_19), .E(n6376), .C(wclk), .QN(n1253) );
  DFE1 \mem_reg_203][18  ( .D(D_18), .E(n6376), .C(wclk), .QN(n1254) );
  DFE1 \mem_reg_203][17  ( .D(D_17), .E(n6376), .C(wclk), .QN(n1255) );
  DFE1 \mem_reg_203][16  ( .D(D_16), .E(n6376), .C(wclk), .QN(n1256) );
  DFE1 \mem_reg_203][15  ( .D(D_15), .E(n6376), .C(wclk), .QN(n1257) );
  DFE1 \mem_reg_203][14  ( .D(D_14), .E(n6376), .C(wclk), .QN(n1258) );
  DFE1 \mem_reg_203][13  ( .D(D_13), .E(n6376), .C(wclk), .QN(n1259) );
  DFE1 \mem_reg_203][12  ( .D(D_12), .E(n6376), .C(wclk), .QN(n1260) );
  DFE1 \mem_reg_203][11  ( .D(D_11), .E(n6376), .C(wclk), .QN(n1261) );
  DFE1 \mem_reg_203][10  ( .D(D_10), .E(n6376), .C(wclk), .QN(n1262) );
  DFE1 \mem_reg_203][9  ( .D(D_9), .E(n6376), .C(wclk), .QN(n1263) );
  DFE1 \mem_reg_203][8  ( .D(D_8), .E(n6376), .C(wclk), .QN(n1264) );
  DFE1 \mem_reg_203][7  ( .D(D_7), .E(n6376), .C(wclk), .QN(n1265) );
  DFE1 \mem_reg_203][6  ( .D(D_6), .E(n6376), .C(wclk), .QN(n1266) );
  DFE1 \mem_reg_203][5  ( .D(D_5), .E(n6376), .C(wclk), .QN(n1267) );
  DFE1 \mem_reg_203][4  ( .D(D_4), .E(n6376), .C(wclk), .QN(n1268) );
  DFE1 \mem_reg_203][3  ( .D(D_3), .E(n6376), .C(wclk), .QN(n1269) );
  DFE1 \mem_reg_203][2  ( .D(D_2), .E(n6376), .C(wclk), .QN(n1270) );
  DFE1 \mem_reg_203][1  ( .D(D_1), .E(n6376), .C(wclk), .QN(n1271) );
  DFE1 \mem_reg_203][0  ( .D(D_0), .E(n6376), .C(wclk), .QN(n1272) );
  DFE1 \mem_reg_202][23  ( .D(D_23), .E(n6375), .C(wclk), .QN(n1273) );
  DFE1 \mem_reg_202][22  ( .D(D_22), .E(n6375), .C(wclk), .QN(n1274) );
  DFE1 \mem_reg_202][21  ( .D(D_21), .E(n6375), .C(wclk), .QN(n1275) );
  DFE1 \mem_reg_202][20  ( .D(D_20), .E(n6375), .C(wclk), .QN(n1276) );
  DFE1 \mem_reg_202][19  ( .D(D_19), .E(n6375), .C(wclk), .QN(n1277) );
  DFE1 \mem_reg_202][18  ( .D(D_18), .E(n6375), .C(wclk), .QN(n1278) );
  DFE1 \mem_reg_202][17  ( .D(D_17), .E(n6375), .C(wclk), .QN(n1279) );
  DFE1 \mem_reg_202][16  ( .D(D_16), .E(n6375), .C(wclk), .QN(n1280) );
  DFE1 \mem_reg_202][15  ( .D(D_15), .E(n6375), .C(wclk), .QN(n1281) );
  DFE1 \mem_reg_202][14  ( .D(D_14), .E(n6375), .C(wclk), .QN(n1282) );
  DFE1 \mem_reg_202][13  ( .D(D_13), .E(n6375), .C(wclk), .QN(n1283) );
  DFE1 \mem_reg_202][12  ( .D(D_12), .E(n6375), .C(wclk), .QN(n1284) );
  DFE1 \mem_reg_202][11  ( .D(D_11), .E(n6375), .C(wclk), .QN(n1285) );
  DFE1 \mem_reg_202][10  ( .D(D_10), .E(n6375), .C(wclk), .QN(n1286) );
  DFE1 \mem_reg_202][9  ( .D(D_9), .E(n6375), .C(wclk), .QN(n1287) );
  DFE1 \mem_reg_202][8  ( .D(D_8), .E(n6375), .C(wclk), .QN(n1288) );
  DFE1 \mem_reg_202][7  ( .D(D_7), .E(n6375), .C(wclk), .QN(n1289) );
  DFE1 \mem_reg_202][6  ( .D(D_6), .E(n6375), .C(wclk), .QN(n1290) );
  DFE1 \mem_reg_202][5  ( .D(D_5), .E(n6375), .C(wclk), .QN(n1291) );
  DFE1 \mem_reg_202][4  ( .D(D_4), .E(n6375), .C(wclk), .QN(n1292) );
  DFE1 \mem_reg_202][3  ( .D(D_3), .E(n6375), .C(wclk), .QN(n1293) );
  DFE1 \mem_reg_202][2  ( .D(D_2), .E(n6375), .C(wclk), .QN(n1294) );
  DFE1 \mem_reg_202][1  ( .D(D_1), .E(n6375), .C(wclk), .QN(n1295) );
  DFE1 \mem_reg_202][0  ( .D(D_0), .E(n6375), .C(wclk), .QN(n1296) );
  DFE1 \mem_reg_201][23  ( .D(D_23), .E(n6374), .C(wclk), .QN(n1297) );
  DFE1 \mem_reg_201][22  ( .D(D_22), .E(n6374), .C(wclk), .QN(n1298) );
  DFE1 \mem_reg_201][21  ( .D(D_21), .E(n6374), .C(wclk), .QN(n1299) );
  DFE1 \mem_reg_201][20  ( .D(D_20), .E(n6374), .C(wclk), .QN(n1300) );
  DFE1 \mem_reg_201][19  ( .D(D_19), .E(n6374), .C(wclk), .QN(n1301) );
  DFE1 \mem_reg_201][18  ( .D(D_18), .E(n6374), .C(wclk), .QN(n1302) );
  DFE1 \mem_reg_201][17  ( .D(D_17), .E(n6374), .C(wclk), .QN(n1303) );
  DFE1 \mem_reg_201][16  ( .D(D_16), .E(n6374), .C(wclk), .QN(n1304) );
  DFE1 \mem_reg_201][15  ( .D(D_15), .E(n6374), .C(wclk), .QN(n1305) );
  DFE1 \mem_reg_201][14  ( .D(D_14), .E(n6374), .C(wclk), .QN(n1306) );
  DFE1 \mem_reg_201][13  ( .D(D_13), .E(n6374), .C(wclk), .QN(n1307) );
  DFE1 \mem_reg_201][12  ( .D(D_12), .E(n6374), .C(wclk), .QN(n1308) );
  DFE1 \mem_reg_201][11  ( .D(D_11), .E(n6374), .C(wclk), .QN(n1309) );
  DFE1 \mem_reg_201][10  ( .D(D_10), .E(n6374), .C(wclk), .QN(n1310) );
  DFE1 \mem_reg_201][9  ( .D(D_9), .E(n6374), .C(wclk), .QN(n1311) );
  DFE1 \mem_reg_201][8  ( .D(D_8), .E(n6374), .C(wclk), .QN(n1312) );
  DFE1 \mem_reg_201][7  ( .D(D_7), .E(n6374), .C(wclk), .QN(n1313) );
  DFE1 \mem_reg_201][6  ( .D(D_6), .E(n6374), .C(wclk), .QN(n1314) );
  DFE1 \mem_reg_201][5  ( .D(D_5), .E(n6374), .C(wclk), .QN(n1315) );
  DFE1 \mem_reg_201][4  ( .D(D_4), .E(n6374), .C(wclk), .QN(n1316) );
  DFE1 \mem_reg_201][3  ( .D(D_3), .E(n6374), .C(wclk), .QN(n1317) );
  DFE1 \mem_reg_201][2  ( .D(D_2), .E(n6374), .C(wclk), .QN(n1318) );
  DFE1 \mem_reg_201][1  ( .D(D_1), .E(n6374), .C(wclk), .QN(n1319) );
  DFE1 \mem_reg_201][0  ( .D(D_0), .E(n6374), .C(wclk), .QN(n1320) );
  DFE1 \mem_reg_200][23  ( .D(D_23), .E(n6373), .C(wclk), .QN(n1321) );
  DFE1 \mem_reg_200][22  ( .D(D_22), .E(n6373), .C(wclk), .QN(n1322) );
  DFE1 \mem_reg_200][21  ( .D(D_21), .E(n6373), .C(wclk), .QN(n1323) );
  DFE1 \mem_reg_200][20  ( .D(D_20), .E(n6373), .C(wclk), .QN(n1324) );
  DFE1 \mem_reg_200][19  ( .D(D_19), .E(n6373), .C(wclk), .QN(n1325) );
  DFE1 \mem_reg_200][18  ( .D(D_18), .E(n6373), .C(wclk), .QN(n1326) );
  DFE1 \mem_reg_200][17  ( .D(D_17), .E(n6373), .C(wclk), .QN(n1327) );
  DFE1 \mem_reg_200][16  ( .D(D_16), .E(n6373), .C(wclk), .QN(n1328) );
  DFE1 \mem_reg_200][15  ( .D(D_15), .E(n6373), .C(wclk), .QN(n1329) );
  DFE1 \mem_reg_200][14  ( .D(D_14), .E(n6373), .C(wclk), .QN(n1330) );
  DFE1 \mem_reg_200][13  ( .D(D_13), .E(n6373), .C(wclk), .QN(n1331) );
  DFE1 \mem_reg_200][12  ( .D(D_12), .E(n6373), .C(wclk), .QN(n1332) );
  DFE1 \mem_reg_200][11  ( .D(D_11), .E(n6373), .C(wclk), .QN(n1333) );
  DFE1 \mem_reg_200][10  ( .D(D_10), .E(n6373), .C(wclk), .QN(n1334) );
  DFE1 \mem_reg_200][9  ( .D(D_9), .E(n6373), .C(wclk), .QN(n1335) );
  DFE1 \mem_reg_200][8  ( .D(D_8), .E(n6373), .C(wclk), .QN(n1336) );
  DFE1 \mem_reg_200][7  ( .D(D_7), .E(n6373), .C(wclk), .QN(n1337) );
  DFE1 \mem_reg_200][6  ( .D(D_6), .E(n6373), .C(wclk), .QN(n1338) );
  DFE1 \mem_reg_200][5  ( .D(D_5), .E(n6373), .C(wclk), .QN(n1339) );
  DFE1 \mem_reg_200][4  ( .D(D_4), .E(n6373), .C(wclk), .QN(n1340) );
  DFE1 \mem_reg_200][3  ( .D(D_3), .E(n6373), .C(wclk), .QN(n1341) );
  DFE1 \mem_reg_200][2  ( .D(D_2), .E(n6373), .C(wclk), .QN(n1342) );
  DFE1 \mem_reg_200][1  ( .D(D_1), .E(n6373), .C(wclk), .QN(n1343) );
  DFE1 \mem_reg_200][0  ( .D(D_0), .E(n6373), .C(wclk), .QN(n1344) );
  DFE1 \mem_reg_199][23  ( .D(D_23), .E(n6372), .C(wclk), .QN(n1345) );
  DFE1 \mem_reg_199][22  ( .D(D_22), .E(n6372), .C(wclk), .QN(n1346) );
  DFE1 \mem_reg_199][21  ( .D(D_21), .E(n6372), .C(wclk), .QN(n1347) );
  DFE1 \mem_reg_199][20  ( .D(D_20), .E(n6372), .C(wclk), .QN(n1348) );
  DFE1 \mem_reg_199][19  ( .D(D_19), .E(n6372), .C(wclk), .QN(n1349) );
  DFE1 \mem_reg_199][18  ( .D(D_18), .E(n6372), .C(wclk), .QN(n1350) );
  DFE1 \mem_reg_199][17  ( .D(D_17), .E(n6372), .C(wclk), .QN(n1351) );
  DFE1 \mem_reg_199][16  ( .D(D_16), .E(n6372), .C(wclk), .QN(n1352) );
  DFE1 \mem_reg_199][15  ( .D(D_15), .E(n6372), .C(wclk), .QN(n1353) );
  DFE1 \mem_reg_199][14  ( .D(D_14), .E(n6372), .C(wclk), .QN(n1354) );
  DFE1 \mem_reg_199][13  ( .D(D_13), .E(n6372), .C(wclk), .QN(n1355) );
  DFE1 \mem_reg_199][12  ( .D(D_12), .E(n6372), .C(wclk), .QN(n1356) );
  DFE1 \mem_reg_199][11  ( .D(D_11), .E(n6372), .C(wclk), .QN(n1357) );
  DFE1 \mem_reg_199][10  ( .D(D_10), .E(n6372), .C(wclk), .QN(n1358) );
  DFE1 \mem_reg_199][9  ( .D(D_9), .E(n6372), .C(wclk), .QN(n1359) );
  DFE1 \mem_reg_199][8  ( .D(D_8), .E(n6372), .C(wclk), .QN(n1360) );
  DFE1 \mem_reg_199][7  ( .D(D_7), .E(n6372), .C(wclk), .QN(n1361) );
  DFE1 \mem_reg_199][6  ( .D(D_6), .E(n6372), .C(wclk), .QN(n1362) );
  DFE1 \mem_reg_199][5  ( .D(D_5), .E(n6372), .C(wclk), .QN(n1363) );
  DFE1 \mem_reg_199][4  ( .D(D_4), .E(n6372), .C(wclk), .QN(n1364) );
  DFE1 \mem_reg_199][3  ( .D(D_3), .E(n6372), .C(wclk), .QN(n1365) );
  DFE1 \mem_reg_199][2  ( .D(D_2), .E(n6372), .C(wclk), .QN(n1366) );
  DFE1 \mem_reg_199][1  ( .D(D_1), .E(n6372), .C(wclk), .QN(n1367) );
  DFE1 \mem_reg_199][0  ( .D(D_0), .E(n6372), .C(wclk), .QN(n1368) );
  DFE1 \mem_reg_198][23  ( .D(D_23), .E(n6371), .C(wclk), .QN(n1369) );
  DFE1 \mem_reg_198][22  ( .D(D_22), .E(n6371), .C(wclk), .QN(n1370) );
  DFE1 \mem_reg_198][21  ( .D(D_21), .E(n6371), .C(wclk), .QN(n1371) );
  DFE1 \mem_reg_198][20  ( .D(D_20), .E(n6371), .C(wclk), .QN(n1372) );
  DFE1 \mem_reg_198][19  ( .D(D_19), .E(n6371), .C(wclk), .QN(n1373) );
  DFE1 \mem_reg_198][18  ( .D(D_18), .E(n6371), .C(wclk), .QN(n1374) );
  DFE1 \mem_reg_198][17  ( .D(D_17), .E(n6371), .C(wclk), .QN(n1375) );
  DFE1 \mem_reg_198][16  ( .D(D_16), .E(n6371), .C(wclk), .QN(n1376) );
  DFE1 \mem_reg_198][15  ( .D(D_15), .E(n6371), .C(wclk), .QN(n1377) );
  DFE1 \mem_reg_198][14  ( .D(D_14), .E(n6371), .C(wclk), .QN(n1378) );
  DFE1 \mem_reg_198][13  ( .D(D_13), .E(n6371), .C(wclk), .QN(n1379) );
  DFE1 \mem_reg_198][12  ( .D(D_12), .E(n6371), .C(wclk), .QN(n1380) );
  DFE1 \mem_reg_198][11  ( .D(D_11), .E(n6371), .C(wclk), .QN(n1381) );
  DFE1 \mem_reg_198][10  ( .D(D_10), .E(n6371), .C(wclk), .QN(n1382) );
  DFE1 \mem_reg_198][9  ( .D(D_9), .E(n6371), .C(wclk), .QN(n1383) );
  DFE1 \mem_reg_198][8  ( .D(D_8), .E(n6371), .C(wclk), .QN(n1384) );
  DFE1 \mem_reg_198][7  ( .D(D_7), .E(n6371), .C(wclk), .QN(n1385) );
  DFE1 \mem_reg_198][6  ( .D(D_6), .E(n6371), .C(wclk), .QN(n1386) );
  DFE1 \mem_reg_198][5  ( .D(D_5), .E(n6371), .C(wclk), .QN(n1387) );
  DFE1 \mem_reg_198][4  ( .D(D_4), .E(n6371), .C(wclk), .QN(n1388) );
  DFE1 \mem_reg_198][3  ( .D(D_3), .E(n6371), .C(wclk), .QN(n1389) );
  DFE1 \mem_reg_198][2  ( .D(D_2), .E(n6371), .C(wclk), .QN(n1390) );
  DFE1 \mem_reg_198][1  ( .D(D_1), .E(n6371), .C(wclk), .QN(n1391) );
  DFE1 \mem_reg_198][0  ( .D(D_0), .E(n6371), .C(wclk), .QN(n1392) );
  DFE1 \mem_reg_197][23  ( .D(D_23), .E(n6370), .C(wclk), .QN(n1393) );
  DFE1 \mem_reg_197][22  ( .D(D_22), .E(n6370), .C(wclk), .QN(n1394) );
  DFE1 \mem_reg_197][21  ( .D(D_21), .E(n6370), .C(wclk), .QN(n1395) );
  DFE1 \mem_reg_197][20  ( .D(D_20), .E(n6370), .C(wclk), .QN(n1396) );
  DFE1 \mem_reg_197][19  ( .D(D_19), .E(n6370), .C(wclk), .QN(n1397) );
  DFE1 \mem_reg_197][18  ( .D(D_18), .E(n6370), .C(wclk), .QN(n1398) );
  DFE1 \mem_reg_197][17  ( .D(D_17), .E(n6370), .C(wclk), .QN(n1399) );
  DFE1 \mem_reg_197][16  ( .D(D_16), .E(n6370), .C(wclk), .QN(n1400) );
  DFE1 \mem_reg_197][15  ( .D(D_15), .E(n6370), .C(wclk), .QN(n1401) );
  DFE1 \mem_reg_197][14  ( .D(D_14), .E(n6370), .C(wclk), .QN(n1402) );
  DFE1 \mem_reg_197][13  ( .D(D_13), .E(n6370), .C(wclk), .QN(n1403) );
  DFE1 \mem_reg_197][12  ( .D(D_12), .E(n6370), .C(wclk), .QN(n1404) );
  DFE1 \mem_reg_197][11  ( .D(D_11), .E(n6370), .C(wclk), .QN(n1405) );
  DFE1 \mem_reg_197][10  ( .D(D_10), .E(n6370), .C(wclk), .QN(n1406) );
  DFE1 \mem_reg_197][9  ( .D(D_9), .E(n6370), .C(wclk), .QN(n1407) );
  DFE1 \mem_reg_197][8  ( .D(D_8), .E(n6370), .C(wclk), .QN(n1408) );
  DFE1 \mem_reg_197][7  ( .D(D_7), .E(n6370), .C(wclk), .QN(n1409) );
  DFE1 \mem_reg_197][6  ( .D(D_6), .E(n6370), .C(wclk), .QN(n1410) );
  DFE1 \mem_reg_197][5  ( .D(D_5), .E(n6370), .C(wclk), .QN(n1411) );
  DFE1 \mem_reg_197][4  ( .D(D_4), .E(n6370), .C(wclk), .QN(n1412) );
  DFE1 \mem_reg_197][3  ( .D(D_3), .E(n6370), .C(wclk), .QN(n1413) );
  DFE1 \mem_reg_197][2  ( .D(D_2), .E(n6370), .C(wclk), .QN(n1414) );
  DFE1 \mem_reg_197][1  ( .D(D_1), .E(n6370), .C(wclk), .QN(n1415) );
  DFE1 \mem_reg_197][0  ( .D(D_0), .E(n6370), .C(wclk), .QN(n1416) );
  DFE1 \mem_reg_196][23  ( .D(D_23), .E(n6369), .C(wclk), .QN(n1417) );
  DFE1 \mem_reg_196][22  ( .D(D_22), .E(n6369), .C(wclk), .QN(n1418) );
  DFE1 \mem_reg_196][21  ( .D(D_21), .E(n6369), .C(wclk), .QN(n1419) );
  DFE1 \mem_reg_196][20  ( .D(D_20), .E(n6369), .C(wclk), .QN(n1420) );
  DFE1 \mem_reg_196][19  ( .D(D_19), .E(n6369), .C(wclk), .QN(n1421) );
  DFE1 \mem_reg_196][18  ( .D(D_18), .E(n6369), .C(wclk), .QN(n1422) );
  DFE1 \mem_reg_196][17  ( .D(D_17), .E(n6369), .C(wclk), .QN(n1423) );
  DFE1 \mem_reg_196][16  ( .D(D_16), .E(n6369), .C(wclk), .QN(n1424) );
  DFE1 \mem_reg_196][15  ( .D(D_15), .E(n6369), .C(wclk), .QN(n1425) );
  DFE1 \mem_reg_196][14  ( .D(D_14), .E(n6369), .C(wclk), .QN(n1426) );
  DFE1 \mem_reg_196][13  ( .D(D_13), .E(n6369), .C(wclk), .QN(n1427) );
  DFE1 \mem_reg_196][12  ( .D(D_12), .E(n6369), .C(wclk), .QN(n1428) );
  DFE1 \mem_reg_196][11  ( .D(D_11), .E(n6369), .C(wclk), .QN(n1429) );
  DFE1 \mem_reg_196][10  ( .D(D_10), .E(n6369), .C(wclk), .QN(n1430) );
  DFE1 \mem_reg_196][9  ( .D(D_9), .E(n6369), .C(wclk), .QN(n1431) );
  DFE1 \mem_reg_196][8  ( .D(D_8), .E(n6369), .C(wclk), .QN(n1432) );
  DFE1 \mem_reg_196][7  ( .D(D_7), .E(n6369), .C(wclk), .QN(n1433) );
  DFE1 \mem_reg_196][6  ( .D(D_6), .E(n6369), .C(wclk), .QN(n1434) );
  DFE1 \mem_reg_196][5  ( .D(D_5), .E(n6369), .C(wclk), .QN(n1435) );
  DFE1 \mem_reg_196][4  ( .D(D_4), .E(n6369), .C(wclk), .QN(n1436) );
  DFE1 \mem_reg_196][3  ( .D(D_3), .E(n6369), .C(wclk), .QN(n1437) );
  DFE1 \mem_reg_196][2  ( .D(D_2), .E(n6369), .C(wclk), .QN(n1438) );
  DFE1 \mem_reg_196][1  ( .D(D_1), .E(n6369), .C(wclk), .QN(n1439) );
  DFE1 \mem_reg_196][0  ( .D(D_0), .E(n6369), .C(wclk), .QN(n1440) );
  DFE1 \mem_reg_195][23  ( .D(D_23), .E(n6368), .C(wclk), .QN(n1441) );
  DFE1 \mem_reg_195][22  ( .D(D_22), .E(n6368), .C(wclk), .QN(n1442) );
  DFE1 \mem_reg_195][21  ( .D(D_21), .E(n6368), .C(wclk), .QN(n1443) );
  DFE1 \mem_reg_195][20  ( .D(D_20), .E(n6368), .C(wclk), .QN(n1444) );
  DFE1 \mem_reg_195][19  ( .D(D_19), .E(n6368), .C(wclk), .QN(n1445) );
  DFE1 \mem_reg_195][18  ( .D(D_18), .E(n6368), .C(wclk), .QN(n1446) );
  DFE1 \mem_reg_195][17  ( .D(D_17), .E(n6368), .C(wclk), .QN(n1447) );
  DFE1 \mem_reg_195][16  ( .D(D_16), .E(n6368), .C(wclk), .QN(n1448) );
  DFE1 \mem_reg_195][15  ( .D(D_15), .E(n6368), .C(wclk), .QN(n1449) );
  DFE1 \mem_reg_195][14  ( .D(D_14), .E(n6368), .C(wclk), .QN(n1450) );
  DFE1 \mem_reg_195][13  ( .D(D_13), .E(n6368), .C(wclk), .QN(n1451) );
  DFE1 \mem_reg_195][12  ( .D(D_12), .E(n6368), .C(wclk), .QN(n1452) );
  DFE1 \mem_reg_195][11  ( .D(D_11), .E(n6368), .C(wclk), .QN(n1453) );
  DFE1 \mem_reg_195][10  ( .D(D_10), .E(n6368), .C(wclk), .QN(n1454) );
  DFE1 \mem_reg_195][9  ( .D(D_9), .E(n6368), .C(wclk), .QN(n1455) );
  DFE1 \mem_reg_195][8  ( .D(D_8), .E(n6368), .C(wclk), .QN(n1456) );
  DFE1 \mem_reg_195][7  ( .D(D_7), .E(n6368), .C(wclk), .QN(n1457) );
  DFE1 \mem_reg_195][6  ( .D(D_6), .E(n6368), .C(wclk), .QN(n1458) );
  DFE1 \mem_reg_195][5  ( .D(D_5), .E(n6368), .C(wclk), .QN(n1459) );
  DFE1 \mem_reg_195][4  ( .D(D_4), .E(n6368), .C(wclk), .QN(n1460) );
  DFE1 \mem_reg_195][3  ( .D(D_3), .E(n6368), .C(wclk), .QN(n1461) );
  DFE1 \mem_reg_195][2  ( .D(D_2), .E(n6368), .C(wclk), .QN(n1462) );
  DFE1 \mem_reg_195][1  ( .D(D_1), .E(n6368), .C(wclk), .QN(n1463) );
  DFE1 \mem_reg_195][0  ( .D(D_0), .E(n6368), .C(wclk), .QN(n1464) );
  DFE1 \mem_reg_194][23  ( .D(D_23), .E(n6367), .C(wclk), .QN(n1465) );
  DFE1 \mem_reg_194][22  ( .D(D_22), .E(n6367), .C(wclk), .QN(n1466) );
  DFE1 \mem_reg_194][21  ( .D(D_21), .E(n6367), .C(wclk), .QN(n1467) );
  DFE1 \mem_reg_194][20  ( .D(D_20), .E(n6367), .C(wclk), .QN(n1468) );
  DFE1 \mem_reg_194][19  ( .D(D_19), .E(n6367), .C(wclk), .QN(n1469) );
  DFE1 \mem_reg_194][18  ( .D(D_18), .E(n6367), .C(wclk), .QN(n1470) );
  DFE1 \mem_reg_194][17  ( .D(D_17), .E(n6367), .C(wclk), .QN(n1471) );
  DFE1 \mem_reg_194][16  ( .D(D_16), .E(n6367), .C(wclk), .QN(n1472) );
  DFE1 \mem_reg_194][15  ( .D(D_15), .E(n6367), .C(wclk), .QN(n1473) );
  DFE1 \mem_reg_194][14  ( .D(D_14), .E(n6367), .C(wclk), .QN(n1474) );
  DFE1 \mem_reg_194][13  ( .D(D_13), .E(n6367), .C(wclk), .QN(n1475) );
  DFE1 \mem_reg_194][12  ( .D(D_12), .E(n6367), .C(wclk), .QN(n1476) );
  DFE1 \mem_reg_194][11  ( .D(D_11), .E(n6367), .C(wclk), .QN(n1477) );
  DFE1 \mem_reg_194][10  ( .D(D_10), .E(n6367), .C(wclk), .QN(n1478) );
  DFE1 \mem_reg_194][9  ( .D(D_9), .E(n6367), .C(wclk), .QN(n1479) );
  DFE1 \mem_reg_194][8  ( .D(D_8), .E(n6367), .C(wclk), .QN(n1480) );
  DFE1 \mem_reg_194][7  ( .D(D_7), .E(n6367), .C(wclk), .QN(n1481) );
  DFE1 \mem_reg_194][6  ( .D(D_6), .E(n6367), .C(wclk), .QN(n1482) );
  DFE1 \mem_reg_194][5  ( .D(D_5), .E(n6367), .C(wclk), .QN(n1483) );
  DFE1 \mem_reg_194][4  ( .D(D_4), .E(n6367), .C(wclk), .QN(n1484) );
  DFE1 \mem_reg_194][3  ( .D(D_3), .E(n6367), .C(wclk), .QN(n1485) );
  DFE1 \mem_reg_194][2  ( .D(D_2), .E(n6367), .C(wclk), .QN(n1486) );
  DFE1 \mem_reg_194][1  ( .D(D_1), .E(n6367), .C(wclk), .QN(n1487) );
  DFE1 \mem_reg_194][0  ( .D(D_0), .E(n6367), .C(wclk), .QN(n1488) );
  DFE1 \mem_reg_193][23  ( .D(D_23), .E(n6366), .C(wclk), .QN(n1489) );
  DFE1 \mem_reg_193][22  ( .D(D_22), .E(n6366), .C(wclk), .QN(n1490) );
  DFE1 \mem_reg_193][21  ( .D(D_21), .E(n6366), .C(wclk), .QN(n1491) );
  DFE1 \mem_reg_193][20  ( .D(D_20), .E(n6366), .C(wclk), .QN(n1492) );
  DFE1 \mem_reg_193][19  ( .D(D_19), .E(n6366), .C(wclk), .QN(n1493) );
  DFE1 \mem_reg_193][18  ( .D(D_18), .E(n6366), .C(wclk), .QN(n1494) );
  DFE1 \mem_reg_193][17  ( .D(D_17), .E(n6366), .C(wclk), .QN(n1495) );
  DFE1 \mem_reg_193][16  ( .D(D_16), .E(n6366), .C(wclk), .QN(n1496) );
  DFE1 \mem_reg_193][15  ( .D(D_15), .E(n6366), .C(wclk), .QN(n1497) );
  DFE1 \mem_reg_193][14  ( .D(D_14), .E(n6366), .C(wclk), .QN(n1498) );
  DFE1 \mem_reg_193][13  ( .D(D_13), .E(n6366), .C(wclk), .QN(n1499) );
  DFE1 \mem_reg_193][12  ( .D(D_12), .E(n6366), .C(wclk), .QN(n1500) );
  DFE1 \mem_reg_193][11  ( .D(D_11), .E(n6366), .C(wclk), .QN(n1501) );
  DFE1 \mem_reg_193][10  ( .D(D_10), .E(n6366), .C(wclk), .QN(n1502) );
  DFE1 \mem_reg_193][9  ( .D(D_9), .E(n6366), .C(wclk), .QN(n1503) );
  DFE1 \mem_reg_193][8  ( .D(D_8), .E(n6366), .C(wclk), .QN(n1504) );
  DFE1 \mem_reg_193][7  ( .D(D_7), .E(n6366), .C(wclk), .QN(n1505) );
  DFE1 \mem_reg_193][6  ( .D(D_6), .E(n6366), .C(wclk), .QN(n1506) );
  DFE1 \mem_reg_193][5  ( .D(D_5), .E(n6366), .C(wclk), .QN(n1507) );
  DFE1 \mem_reg_193][4  ( .D(D_4), .E(n6366), .C(wclk), .QN(n1508) );
  DFE1 \mem_reg_193][3  ( .D(D_3), .E(n6366), .C(wclk), .QN(n1509) );
  DFE1 \mem_reg_193][2  ( .D(D_2), .E(n6366), .C(wclk), .QN(n1510) );
  DFE1 \mem_reg_193][1  ( .D(D_1), .E(n6366), .C(wclk), .QN(n1511) );
  DFE1 \mem_reg_193][0  ( .D(D_0), .E(n6366), .C(wclk), .QN(n1512) );
  DFE1 \mem_reg_192][23  ( .D(D_23), .E(n6364), .C(wclk), .QN(n1513) );
  DFE1 \mem_reg_192][22  ( .D(D_22), .E(n6364), .C(wclk), .QN(n1514) );
  DFE1 \mem_reg_192][21  ( .D(D_21), .E(n6364), .C(wclk), .QN(n1515) );
  DFE1 \mem_reg_192][20  ( .D(D_20), .E(n6364), .C(wclk), .QN(n1516) );
  DFE1 \mem_reg_192][19  ( .D(D_19), .E(n6364), .C(wclk), .QN(n1517) );
  DFE1 \mem_reg_192][18  ( .D(D_18), .E(n6364), .C(wclk), .QN(n1518) );
  DFE1 \mem_reg_192][17  ( .D(D_17), .E(n6364), .C(wclk), .QN(n1519) );
  DFE1 \mem_reg_192][16  ( .D(D_16), .E(n6364), .C(wclk), .QN(n1520) );
  DFE1 \mem_reg_192][15  ( .D(D_15), .E(n6364), .C(wclk), .QN(n1521) );
  DFE1 \mem_reg_192][14  ( .D(D_14), .E(n6364), .C(wclk), .QN(n1522) );
  DFE1 \mem_reg_192][13  ( .D(D_13), .E(n6364), .C(wclk), .QN(n1523) );
  DFE1 \mem_reg_192][12  ( .D(D_12), .E(n6364), .C(wclk), .QN(n1524) );
  DFE1 \mem_reg_192][11  ( .D(D_11), .E(n6364), .C(wclk), .QN(n1525) );
  DFE1 \mem_reg_192][10  ( .D(D_10), .E(n6364), .C(wclk), .QN(n1526) );
  DFE1 \mem_reg_192][9  ( .D(D_9), .E(n6364), .C(wclk), .QN(n1527) );
  DFE1 \mem_reg_192][8  ( .D(D_8), .E(n6364), .C(wclk), .QN(n1528) );
  DFE1 \mem_reg_192][7  ( .D(D_7), .E(n6364), .C(wclk), .QN(n1529) );
  DFE1 \mem_reg_192][6  ( .D(D_6), .E(n6364), .C(wclk), .QN(n1530) );
  DFE1 \mem_reg_192][5  ( .D(D_5), .E(n6364), .C(wclk), .QN(n1531) );
  DFE1 \mem_reg_192][4  ( .D(D_4), .E(n6364), .C(wclk), .QN(n1532) );
  DFE1 \mem_reg_192][3  ( .D(D_3), .E(n6364), .C(wclk), .QN(n1533) );
  DFE1 \mem_reg_192][2  ( .D(D_2), .E(n6364), .C(wclk), .QN(n1534) );
  DFE1 \mem_reg_192][1  ( .D(D_1), .E(n6364), .C(wclk), .QN(n1535) );
  DFE1 \mem_reg_192][0  ( .D(D_0), .E(n6364), .C(wclk), .QN(n1536) );
  DFE1 \mem_reg_59][23  ( .D(D_23), .E(n6495), .C(wclk), .QN(n4705) );
  DFE1 \mem_reg_59][22  ( .D(D_22), .E(n6495), .C(wclk), .QN(n4706) );
  DFE1 \mem_reg_59][21  ( .D(D_21), .E(n6495), .C(wclk), .QN(n4707) );
  DFE1 \mem_reg_59][20  ( .D(D_20), .E(n6495), .C(wclk), .QN(n4708) );
  DFE1 \mem_reg_59][19  ( .D(D_19), .E(n6495), .C(wclk), .QN(n4709) );
  DFE1 \mem_reg_59][18  ( .D(D_18), .E(n6495), .C(wclk), .QN(n4710) );
  DFE1 \mem_reg_59][17  ( .D(D_17), .E(n6495), .C(wclk), .QN(n4711) );
  DFE1 \mem_reg_59][16  ( .D(D_16), .E(n6495), .C(wclk), .QN(n4712) );
  DFE1 \mem_reg_59][15  ( .D(D_15), .E(n6495), .C(wclk), .QN(n4713) );
  DFE1 \mem_reg_59][14  ( .D(D_14), .E(n6495), .C(wclk), .QN(n4714) );
  DFE1 \mem_reg_59][13  ( .D(D_13), .E(n6495), .C(wclk), .QN(n4715) );
  DFE1 \mem_reg_59][12  ( .D(D_12), .E(n6495), .C(wclk), .QN(n4716) );
  DFE1 \mem_reg_59][11  ( .D(D_11), .E(n6495), .C(wclk), .QN(n4717) );
  DFE1 \mem_reg_59][10  ( .D(D_10), .E(n6495), .C(wclk), .QN(n4718) );
  DFE1 \mem_reg_59][9  ( .D(D_9), .E(n6495), .C(wclk), .QN(n4719) );
  DFE1 \mem_reg_59][8  ( .D(D_8), .E(n6495), .C(wclk), .QN(n4720) );
  DFE1 \mem_reg_59][7  ( .D(D_7), .E(n6495), .C(wclk), .QN(n4721) );
  DFE1 \mem_reg_59][6  ( .D(D_6), .E(n6495), .C(wclk), .QN(n4722) );
  DFE1 \mem_reg_59][5  ( .D(D_5), .E(n6495), .C(wclk), .QN(n4723) );
  DFE1 \mem_reg_59][4  ( .D(D_4), .E(n6495), .C(wclk), .QN(n4724) );
  DFE1 \mem_reg_59][3  ( .D(D_3), .E(n6495), .C(wclk), .QN(n4725) );
  DFE1 \mem_reg_59][2  ( .D(D_2), .E(n6495), .C(wclk), .QN(n4726) );
  DFE1 \mem_reg_59][1  ( .D(D_1), .E(n6495), .C(wclk), .QN(n4727) );
  DFE1 \mem_reg_59][0  ( .D(D_0), .E(n6495), .C(wclk), .QN(n4728) );
  DFE1 \mem_reg_58][23  ( .D(D_23), .E(n6494), .C(wclk), .QN(n4729) );
  DFE1 \mem_reg_58][22  ( .D(D_22), .E(n6494), .C(wclk), .QN(n4730) );
  DFE1 \mem_reg_58][21  ( .D(D_21), .E(n6494), .C(wclk), .QN(n4731) );
  DFE1 \mem_reg_58][20  ( .D(D_20), .E(n6494), .C(wclk), .QN(n4732) );
  DFE1 \mem_reg_58][19  ( .D(D_19), .E(n6494), .C(wclk), .QN(n4733) );
  DFE1 \mem_reg_58][18  ( .D(D_18), .E(n6494), .C(wclk), .QN(n4734) );
  DFE1 \mem_reg_58][17  ( .D(D_17), .E(n6494), .C(wclk), .QN(n4735) );
  DFE1 \mem_reg_58][16  ( .D(D_16), .E(n6494), .C(wclk), .QN(n4736) );
  DFE1 \mem_reg_58][15  ( .D(D_15), .E(n6494), .C(wclk), .QN(n4737) );
  DFE1 \mem_reg_58][14  ( .D(D_14), .E(n6494), .C(wclk), .QN(n4738) );
  DFE1 \mem_reg_58][13  ( .D(D_13), .E(n6494), .C(wclk), .QN(n4739) );
  DFE1 \mem_reg_58][12  ( .D(D_12), .E(n6494), .C(wclk), .QN(n4740) );
  DFE1 \mem_reg_58][11  ( .D(D_11), .E(n6494), .C(wclk), .QN(n4741) );
  DFE1 \mem_reg_58][10  ( .D(D_10), .E(n6494), .C(wclk), .QN(n4742) );
  DFE1 \mem_reg_58][9  ( .D(D_9), .E(n6494), .C(wclk), .QN(n4743) );
  DFE1 \mem_reg_58][8  ( .D(D_8), .E(n6494), .C(wclk), .QN(n4744) );
  DFE1 \mem_reg_58][7  ( .D(D_7), .E(n6494), .C(wclk), .QN(n4745) );
  DFE1 \mem_reg_58][6  ( .D(D_6), .E(n6494), .C(wclk), .QN(n4746) );
  DFE1 \mem_reg_58][5  ( .D(D_5), .E(n6494), .C(wclk), .QN(n4747) );
  DFE1 \mem_reg_58][4  ( .D(D_4), .E(n6494), .C(wclk), .QN(n4748) );
  DFE1 \mem_reg_58][3  ( .D(D_3), .E(n6494), .C(wclk), .QN(n4749) );
  DFE1 \mem_reg_58][2  ( .D(D_2), .E(n6494), .C(wclk), .QN(n4750) );
  DFE1 \mem_reg_58][1  ( .D(D_1), .E(n6494), .C(wclk), .QN(n4751) );
  DFE1 \mem_reg_58][0  ( .D(D_0), .E(n6494), .C(wclk), .QN(n4752) );
  DFE1 \mem_reg_61][23  ( .D(D_23), .E(n6193), .C(wclk), .QN(n4657) );
  DFE1 \mem_reg_61][22  ( .D(D_22), .E(n6193), .C(wclk), .QN(n4658) );
  DFE1 \mem_reg_61][21  ( .D(D_21), .E(n6193), .C(wclk), .QN(n4659) );
  DFE1 \mem_reg_61][20  ( .D(D_20), .E(n6193), .C(wclk), .QN(n4660) );
  DFE1 \mem_reg_61][19  ( .D(D_19), .E(n6193), .C(wclk), .QN(n4661) );
  DFE1 \mem_reg_61][18  ( .D(D_18), .E(n6193), .C(wclk), .QN(n4662) );
  DFE1 \mem_reg_61][17  ( .D(D_17), .E(n6193), .C(wclk), .QN(n4663) );
  DFE1 \mem_reg_61][16  ( .D(D_16), .E(n6193), .C(wclk), .QN(n4664) );
  DFE1 \mem_reg_61][15  ( .D(D_15), .E(n6193), .C(wclk), .QN(n4665) );
  DFE1 \mem_reg_61][14  ( .D(D_14), .E(n6193), .C(wclk), .QN(n4666) );
  DFE1 \mem_reg_61][13  ( .D(D_13), .E(n6193), .C(wclk), .QN(n4667) );
  DFE1 \mem_reg_61][12  ( .D(D_12), .E(n6193), .C(wclk), .QN(n4668) );
  DFE1 \mem_reg_61][11  ( .D(D_11), .E(n6193), .C(wclk), .QN(n4669) );
  DFE1 \mem_reg_61][10  ( .D(D_10), .E(n6193), .C(wclk), .QN(n4670) );
  DFE1 \mem_reg_61][9  ( .D(D_9), .E(n6193), .C(wclk), .QN(n4671) );
  DFE1 \mem_reg_61][8  ( .D(D_8), .E(n6193), .C(wclk), .QN(n4672) );
  DFE1 \mem_reg_61][7  ( .D(D_7), .E(n6193), .C(wclk), .QN(n4673) );
  DFE1 \mem_reg_61][6  ( .D(D_6), .E(n6193), .C(wclk), .QN(n4674) );
  DFE1 \mem_reg_61][5  ( .D(D_5), .E(n6193), .C(wclk), .QN(n4675) );
  DFE1 \mem_reg_61][4  ( .D(D_4), .E(n6193), .C(wclk), .QN(n4676) );
  DFE1 \mem_reg_61][3  ( .D(D_3), .E(n6193), .C(wclk), .QN(n4677) );
  DFE1 \mem_reg_61][2  ( .D(D_2), .E(n6193), .C(wclk), .QN(n4678) );
  DFE1 \mem_reg_61][1  ( .D(D_1), .E(n6193), .C(wclk), .QN(n4679) );
  DFE1 \mem_reg_61][0  ( .D(D_0), .E(n6193), .C(wclk), .QN(n4680) );
  DFE1 \mem_reg_247][23  ( .D(D_23), .E(n6471), .C(wclk), .QN(n193) );
  DFE1 \mem_reg_247][22  ( .D(D_22), .E(n6471), .C(wclk), .QN(n194) );
  DFE1 \mem_reg_247][21  ( .D(D_21), .E(n6471), .C(wclk), .QN(n195) );
  DFE1 \mem_reg_247][20  ( .D(D_20), .E(n6471), .C(wclk), .QN(n196) );
  DFE1 \mem_reg_247][19  ( .D(D_19), .E(n6471), .C(wclk), .QN(n197) );
  DFE1 \mem_reg_247][18  ( .D(D_18), .E(n6471), .C(wclk), .QN(n198) );
  DFE1 \mem_reg_247][17  ( .D(D_17), .E(n6471), .C(wclk), .QN(n199) );
  DFE1 \mem_reg_247][16  ( .D(D_16), .E(n6471), .C(wclk), .QN(n200) );
  DFE1 \mem_reg_247][15  ( .D(D_15), .E(n6471), .C(wclk), .QN(n201) );
  DFE1 \mem_reg_247][14  ( .D(D_14), .E(n6471), .C(wclk), .QN(n202) );
  DFE1 \mem_reg_247][13  ( .D(D_13), .E(n6471), .C(wclk), .QN(n203) );
  DFE1 \mem_reg_247][12  ( .D(D_12), .E(n6471), .C(wclk), .QN(n204) );
  DFE1 \mem_reg_247][11  ( .D(D_11), .E(n6471), .C(wclk), .QN(n205) );
  DFE1 \mem_reg_247][10  ( .D(D_10), .E(n6471), .C(wclk), .QN(n206) );
  DFE1 \mem_reg_247][9  ( .D(D_9), .E(n6471), .C(wclk), .QN(n207) );
  DFE1 \mem_reg_247][8  ( .D(D_8), .E(n6471), .C(wclk), .QN(n208) );
  DFE1 \mem_reg_247][7  ( .D(D_7), .E(n6471), .C(wclk), .QN(n209) );
  DFE1 \mem_reg_247][6  ( .D(D_6), .E(n6471), .C(wclk), .QN(n210) );
  DFE1 \mem_reg_247][5  ( .D(D_5), .E(n6471), .C(wclk), .QN(n211) );
  DFE1 \mem_reg_247][4  ( .D(D_4), .E(n6471), .C(wclk), .QN(n212) );
  DFE1 \mem_reg_247][3  ( .D(D_3), .E(n6471), .C(wclk), .QN(n213) );
  DFE1 \mem_reg_247][2  ( .D(D_2), .E(n6471), .C(wclk), .QN(n214) );
  DFE1 \mem_reg_247][1  ( .D(D_1), .E(n6471), .C(wclk), .QN(n215) );
  DFE1 \mem_reg_247][0  ( .D(D_0), .E(n6471), .C(wclk), .QN(n216) );
  DFE1 \mem_reg_246][23  ( .D(D_23), .E(n6460), .C(wclk), .QN(n217) );
  DFE1 \mem_reg_246][22  ( .D(D_22), .E(n6460), .C(wclk), .QN(n218) );
  DFE1 \mem_reg_246][21  ( .D(D_21), .E(n6460), .C(wclk), .QN(n219) );
  DFE1 \mem_reg_246][20  ( .D(D_20), .E(n6460), .C(wclk), .QN(n220) );
  DFE1 \mem_reg_246][19  ( .D(D_19), .E(n6460), .C(wclk), .QN(n221) );
  DFE1 \mem_reg_246][18  ( .D(D_18), .E(n6460), .C(wclk), .QN(n222) );
  DFE1 \mem_reg_246][17  ( .D(D_17), .E(n6460), .C(wclk), .QN(n223) );
  DFE1 \mem_reg_246][16  ( .D(D_16), .E(n6460), .C(wclk), .QN(n224) );
  DFE1 \mem_reg_246][15  ( .D(D_15), .E(n6460), .C(wclk), .QN(n225) );
  DFE1 \mem_reg_246][14  ( .D(D_14), .E(n6460), .C(wclk), .QN(n226) );
  DFE1 \mem_reg_246][13  ( .D(D_13), .E(n6460), .C(wclk), .QN(n227) );
  DFE1 \mem_reg_246][12  ( .D(D_12), .E(n6460), .C(wclk), .QN(n228) );
  DFE1 \mem_reg_246][11  ( .D(D_11), .E(n6460), .C(wclk), .QN(n229) );
  DFE1 \mem_reg_246][10  ( .D(D_10), .E(n6460), .C(wclk), .QN(n230) );
  DFE1 \mem_reg_246][9  ( .D(D_9), .E(n6460), .C(wclk), .QN(n231) );
  DFE1 \mem_reg_246][8  ( .D(D_8), .E(n6460), .C(wclk), .QN(n232) );
  DFE1 \mem_reg_246][7  ( .D(D_7), .E(n6460), .C(wclk), .QN(n233) );
  DFE1 \mem_reg_246][6  ( .D(D_6), .E(n6460), .C(wclk), .QN(n234) );
  DFE1 \mem_reg_246][5  ( .D(D_5), .E(n6460), .C(wclk), .QN(n235) );
  DFE1 \mem_reg_246][4  ( .D(D_4), .E(n6460), .C(wclk), .QN(n236) );
  DFE1 \mem_reg_246][3  ( .D(D_3), .E(n6460), .C(wclk), .QN(n237) );
  DFE1 \mem_reg_246][2  ( .D(D_2), .E(n6460), .C(wclk), .QN(n238) );
  DFE1 \mem_reg_246][1  ( .D(D_1), .E(n6460), .C(wclk), .QN(n239) );
  DFE1 \mem_reg_246][0  ( .D(D_0), .E(n6460), .C(wclk), .QN(n240) );
  DFE1 \mem_reg_243][23  ( .D(D_23), .E(n6424), .C(wclk), .QN(n289) );
  DFE1 \mem_reg_243][22  ( .D(D_22), .E(n6424), .C(wclk), .QN(n290) );
  DFE1 \mem_reg_243][21  ( .D(D_21), .E(n6424), .C(wclk), .QN(n291) );
  DFE1 \mem_reg_243][20  ( .D(D_20), .E(n6424), .C(wclk), .QN(n292) );
  DFE1 \mem_reg_243][19  ( .D(D_19), .E(n6424), .C(wclk), .QN(n293) );
  DFE1 \mem_reg_243][18  ( .D(D_18), .E(n6424), .C(wclk), .QN(n294) );
  DFE1 \mem_reg_243][17  ( .D(D_17), .E(n6424), .C(wclk), .QN(n295) );
  DFE1 \mem_reg_243][16  ( .D(D_16), .E(n6424), .C(wclk), .QN(n296) );
  DFE1 \mem_reg_243][15  ( .D(D_15), .E(n6424), .C(wclk), .QN(n297) );
  DFE1 \mem_reg_243][14  ( .D(D_14), .E(n6424), .C(wclk), .QN(n298) );
  DFE1 \mem_reg_243][13  ( .D(D_13), .E(n6424), .C(wclk), .QN(n299) );
  DFE1 \mem_reg_243][12  ( .D(D_12), .E(n6424), .C(wclk), .QN(n300) );
  DFE1 \mem_reg_243][11  ( .D(D_11), .E(n6424), .C(wclk), .QN(n301) );
  DFE1 \mem_reg_243][10  ( .D(D_10), .E(n6424), .C(wclk), .QN(n302) );
  DFE1 \mem_reg_243][9  ( .D(D_9), .E(n6424), .C(wclk), .QN(n303) );
  DFE1 \mem_reg_243][8  ( .D(D_8), .E(n6424), .C(wclk), .QN(n304) );
  DFE1 \mem_reg_243][7  ( .D(D_7), .E(n6424), .C(wclk), .QN(n305) );
  DFE1 \mem_reg_243][6  ( .D(D_6), .E(n6424), .C(wclk), .QN(n306) );
  DFE1 \mem_reg_243][5  ( .D(D_5), .E(n6424), .C(wclk), .QN(n307) );
  DFE1 \mem_reg_243][4  ( .D(D_4), .E(n6424), .C(wclk), .QN(n308) );
  DFE1 \mem_reg_243][3  ( .D(D_3), .E(n6424), .C(wclk), .QN(n309) );
  DFE1 \mem_reg_243][2  ( .D(D_2), .E(n6424), .C(wclk), .QN(n310) );
  DFE1 \mem_reg_243][1  ( .D(D_1), .E(n6424), .C(wclk), .QN(n311) );
  DFE1 \mem_reg_243][0  ( .D(D_0), .E(n6424), .C(wclk), .QN(n312) );
  DFE1 \mem_reg_242][23  ( .D(D_23), .E(n6418), .C(wclk), .QN(n313) );
  DFE1 \mem_reg_242][22  ( .D(D_22), .E(n6418), .C(wclk), .QN(n314) );
  DFE1 \mem_reg_242][21  ( .D(D_21), .E(n6418), .C(wclk), .QN(n315) );
  DFE1 \mem_reg_242][20  ( .D(D_20), .E(n6418), .C(wclk), .QN(n316) );
  DFE1 \mem_reg_242][19  ( .D(D_19), .E(n6418), .C(wclk), .QN(n317) );
  DFE1 \mem_reg_242][18  ( .D(D_18), .E(n6418), .C(wclk), .QN(n318) );
  DFE1 \mem_reg_242][17  ( .D(D_17), .E(n6418), .C(wclk), .QN(n319) );
  DFE1 \mem_reg_242][16  ( .D(D_16), .E(n6418), .C(wclk), .QN(n320) );
  DFE1 \mem_reg_242][15  ( .D(D_15), .E(n6418), .C(wclk), .QN(n321) );
  DFE1 \mem_reg_242][14  ( .D(D_14), .E(n6418), .C(wclk), .QN(n322) );
  DFE1 \mem_reg_242][13  ( .D(D_13), .E(n6418), .C(wclk), .QN(n323) );
  DFE1 \mem_reg_242][12  ( .D(D_12), .E(n6418), .C(wclk), .QN(n324) );
  DFE1 \mem_reg_242][11  ( .D(D_11), .E(n6418), .C(wclk), .QN(n325) );
  DFE1 \mem_reg_242][10  ( .D(D_10), .E(n6418), .C(wclk), .QN(n326) );
  DFE1 \mem_reg_242][9  ( .D(D_9), .E(n6418), .C(wclk), .QN(n327) );
  DFE1 \mem_reg_242][8  ( .D(D_8), .E(n6418), .C(wclk), .QN(n328) );
  DFE1 \mem_reg_242][7  ( .D(D_7), .E(n6418), .C(wclk), .QN(n329) );
  DFE1 \mem_reg_242][6  ( .D(D_6), .E(n6418), .C(wclk), .QN(n330) );
  DFE1 \mem_reg_242][5  ( .D(D_5), .E(n6418), .C(wclk), .QN(n331) );
  DFE1 \mem_reg_242][4  ( .D(D_4), .E(n6418), .C(wclk), .QN(n332) );
  DFE1 \mem_reg_242][3  ( .D(D_3), .E(n6418), .C(wclk), .QN(n333) );
  DFE1 \mem_reg_242][2  ( .D(D_2), .E(n6418), .C(wclk), .QN(n334) );
  DFE1 \mem_reg_242][1  ( .D(D_1), .E(n6418), .C(wclk), .QN(n335) );
  DFE1 \mem_reg_242][0  ( .D(D_0), .E(n6418), .C(wclk), .QN(n336) );
  DFE1 \mem_reg_255][23  ( .D(D_23), .E(n6289), .C(wclk), .QN(n1) );
  DFE1 \mem_reg_255][22  ( .D(D_22), .E(n6289), .C(wclk), .QN(n2) );
  DFE1 \mem_reg_255][21  ( .D(D_21), .E(n6289), .C(wclk), .QN(n3) );
  DFE1 \mem_reg_255][20  ( .D(D_20), .E(n6289), .C(wclk), .QN(n4) );
  DFE1 \mem_reg_255][19  ( .D(D_19), .E(n6289), .C(wclk), .QN(n5) );
  DFE1 \mem_reg_255][18  ( .D(D_18), .E(n6289), .C(wclk), .QN(n6) );
  DFE1 \mem_reg_255][17  ( .D(D_17), .E(n6289), .C(wclk), .QN(n7) );
  DFE1 \mem_reg_255][16  ( .D(D_16), .E(n6289), .C(wclk), .QN(n8) );
  DFE1 \mem_reg_255][15  ( .D(D_15), .E(n6289), .C(wclk), .QN(n9) );
  DFE1 \mem_reg_255][14  ( .D(D_14), .E(n6289), .C(wclk), .QN(n10) );
  DFE1 \mem_reg_255][13  ( .D(D_13), .E(n6289), .C(wclk), .QN(n11) );
  DFE1 \mem_reg_255][12  ( .D(D_12), .E(n6289), .C(wclk), .QN(n12) );
  DFE1 \mem_reg_255][11  ( .D(D_11), .E(n6289), .C(wclk), .QN(n13) );
  DFE1 \mem_reg_255][10  ( .D(D_10), .E(n6289), .C(wclk), .QN(n14) );
  DFE1 \mem_reg_255][9  ( .D(D_9), .E(n6289), .C(wclk), .QN(n15) );
  DFE1 \mem_reg_255][8  ( .D(D_8), .E(n6289), .C(wclk), .QN(n16) );
  DFE1 \mem_reg_255][7  ( .D(D_7), .E(n6289), .C(wclk), .QN(n17) );
  DFE1 \mem_reg_255][6  ( .D(D_6), .E(n6289), .C(wclk), .QN(n18) );
  DFE1 \mem_reg_255][5  ( .D(D_5), .E(n6289), .C(wclk), .QN(n19) );
  DFE1 \mem_reg_255][4  ( .D(D_4), .E(n6289), .C(wclk), .QN(n20) );
  DFE1 \mem_reg_255][3  ( .D(D_3), .E(n6289), .C(wclk), .QN(n21) );
  DFE1 \mem_reg_255][2  ( .D(D_2), .E(n6289), .C(wclk), .QN(n22) );
  DFE1 \mem_reg_255][1  ( .D(D_1), .E(n6289), .C(wclk), .QN(n23) );
  DFE1 \mem_reg_255][0  ( .D(D_0), .E(n6289), .C(wclk), .QN(n24) );
  DFE1 \mem_reg_254][23  ( .D(D_23), .E(n6278), .C(wclk), .QN(n25) );
  DFE1 \mem_reg_254][22  ( .D(D_22), .E(n6278), .C(wclk), .QN(n26) );
  DFE1 \mem_reg_254][21  ( .D(D_21), .E(n6278), .C(wclk), .QN(n27) );
  DFE1 \mem_reg_254][20  ( .D(D_20), .E(n6278), .C(wclk), .QN(n28) );
  DFE1 \mem_reg_254][19  ( .D(D_19), .E(n6278), .C(wclk), .QN(n29) );
  DFE1 \mem_reg_254][18  ( .D(D_18), .E(n6278), .C(wclk), .QN(n30) );
  DFE1 \mem_reg_254][17  ( .D(D_17), .E(n6278), .C(wclk), .QN(n31) );
  DFE1 \mem_reg_254][16  ( .D(D_16), .E(n6278), .C(wclk), .QN(n32) );
  DFE1 \mem_reg_254][15  ( .D(D_15), .E(n6278), .C(wclk), .QN(n33) );
  DFE1 \mem_reg_254][14  ( .D(D_14), .E(n6278), .C(wclk), .QN(n34) );
  DFE1 \mem_reg_254][13  ( .D(D_13), .E(n6278), .C(wclk), .QN(n35) );
  DFE1 \mem_reg_254][12  ( .D(D_12), .E(n6278), .C(wclk), .QN(n36) );
  DFE1 \mem_reg_254][11  ( .D(D_11), .E(n6278), .C(wclk), .QN(n37) );
  DFE1 \mem_reg_254][10  ( .D(D_10), .E(n6278), .C(wclk), .QN(n38) );
  DFE1 \mem_reg_254][9  ( .D(D_9), .E(n6278), .C(wclk), .QN(n39) );
  DFE1 \mem_reg_254][8  ( .D(D_8), .E(n6278), .C(wclk), .QN(n40) );
  DFE1 \mem_reg_254][7  ( .D(D_7), .E(n6278), .C(wclk), .QN(n41) );
  DFE1 \mem_reg_254][6  ( .D(D_6), .E(n6278), .C(wclk), .QN(n42) );
  DFE1 \mem_reg_254][5  ( .D(D_5), .E(n6278), .C(wclk), .QN(n43) );
  DFE1 \mem_reg_254][4  ( .D(D_4), .E(n6278), .C(wclk), .QN(n44) );
  DFE1 \mem_reg_254][3  ( .D(D_3), .E(n6278), .C(wclk), .QN(n45) );
  DFE1 \mem_reg_254][2  ( .D(D_2), .E(n6278), .C(wclk), .QN(n46) );
  DFE1 \mem_reg_254][1  ( .D(D_1), .E(n6278), .C(wclk), .QN(n47) );
  DFE1 \mem_reg_254][0  ( .D(D_0), .E(n6278), .C(wclk), .QN(n48) );
  DFE1 \mem_reg_252][23  ( .D(D_23), .E(n6252), .C(wclk), .QN(n73) );
  DFE1 \mem_reg_252][22  ( .D(D_22), .E(n6252), .C(wclk), .QN(n74) );
  DFE1 \mem_reg_252][21  ( .D(D_21), .E(n6252), .C(wclk), .QN(n75) );
  DFE1 \mem_reg_252][20  ( .D(D_20), .E(n6252), .C(wclk), .QN(n76) );
  DFE1 \mem_reg_252][19  ( .D(D_19), .E(n6252), .C(wclk), .QN(n77) );
  DFE1 \mem_reg_252][18  ( .D(D_18), .E(n6252), .C(wclk), .QN(n78) );
  DFE1 \mem_reg_252][17  ( .D(D_17), .E(n6252), .C(wclk), .QN(n79) );
  DFE1 \mem_reg_252][16  ( .D(D_16), .E(n6252), .C(wclk), .QN(n80) );
  DFE1 \mem_reg_252][15  ( .D(D_15), .E(n6252), .C(wclk), .QN(n81) );
  DFE1 \mem_reg_252][14  ( .D(D_14), .E(n6252), .C(wclk), .QN(n82) );
  DFE1 \mem_reg_252][13  ( .D(D_13), .E(n6252), .C(wclk), .QN(n83) );
  DFE1 \mem_reg_252][12  ( .D(D_12), .E(n6252), .C(wclk), .QN(n84) );
  DFE1 \mem_reg_252][11  ( .D(D_11), .E(n6252), .C(wclk), .QN(n85) );
  DFE1 \mem_reg_252][10  ( .D(D_10), .E(n6252), .C(wclk), .QN(n86) );
  DFE1 \mem_reg_252][9  ( .D(D_9), .E(n6252), .C(wclk), .QN(n87) );
  DFE1 \mem_reg_252][8  ( .D(D_8), .E(n6252), .C(wclk), .QN(n88) );
  DFE1 \mem_reg_252][7  ( .D(D_7), .E(n6252), .C(wclk), .QN(n89) );
  DFE1 \mem_reg_252][6  ( .D(D_6), .E(n6252), .C(wclk), .QN(n90) );
  DFE1 \mem_reg_252][5  ( .D(D_5), .E(n6252), .C(wclk), .QN(n91) );
  DFE1 \mem_reg_252][4  ( .D(D_4), .E(n6252), .C(wclk), .QN(n92) );
  DFE1 \mem_reg_252][3  ( .D(D_3), .E(n6252), .C(wclk), .QN(n93) );
  DFE1 \mem_reg_252][2  ( .D(D_2), .E(n6252), .C(wclk), .QN(n94) );
  DFE1 \mem_reg_252][1  ( .D(D_1), .E(n6252), .C(wclk), .QN(n95) );
  DFE1 \mem_reg_252][0  ( .D(D_0), .E(n6252), .C(wclk), .QN(n96) );
  DFE1 \mem_reg_244][23  ( .D(D_23), .E(n6435), .C(wclk), .QN(n265) );
  DFE1 \mem_reg_244][22  ( .D(D_22), .E(n6435), .C(wclk), .QN(n266) );
  DFE1 \mem_reg_244][21  ( .D(D_21), .E(n6435), .C(wclk), .QN(n267) );
  DFE1 \mem_reg_244][20  ( .D(D_20), .E(n6435), .C(wclk), .QN(n268) );
  DFE1 \mem_reg_244][19  ( .D(D_19), .E(n6435), .C(wclk), .QN(n269) );
  DFE1 \mem_reg_244][18  ( .D(D_18), .E(n6435), .C(wclk), .QN(n270) );
  DFE1 \mem_reg_244][17  ( .D(D_17), .E(n6435), .C(wclk), .QN(n271) );
  DFE1 \mem_reg_244][16  ( .D(D_16), .E(n6435), .C(wclk), .QN(n272) );
  DFE1 \mem_reg_244][15  ( .D(D_15), .E(n6435), .C(wclk), .QN(n273) );
  DFE1 \mem_reg_244][14  ( .D(D_14), .E(n6435), .C(wclk), .QN(n274) );
  DFE1 \mem_reg_244][13  ( .D(D_13), .E(n6435), .C(wclk), .QN(n275) );
  DFE1 \mem_reg_244][12  ( .D(D_12), .E(n6435), .C(wclk), .QN(n276) );
  DFE1 \mem_reg_244][11  ( .D(D_11), .E(n6435), .C(wclk), .QN(n277) );
  DFE1 \mem_reg_244][10  ( .D(D_10), .E(n6435), .C(wclk), .QN(n278) );
  DFE1 \mem_reg_244][9  ( .D(D_9), .E(n6435), .C(wclk), .QN(n279) );
  DFE1 \mem_reg_244][8  ( .D(D_8), .E(n6435), .C(wclk), .QN(n280) );
  DFE1 \mem_reg_244][7  ( .D(D_7), .E(n6435), .C(wclk), .QN(n281) );
  DFE1 \mem_reg_244][6  ( .D(D_6), .E(n6435), .C(wclk), .QN(n282) );
  DFE1 \mem_reg_244][5  ( .D(D_5), .E(n6435), .C(wclk), .QN(n283) );
  DFE1 \mem_reg_244][4  ( .D(D_4), .E(n6435), .C(wclk), .QN(n284) );
  DFE1 \mem_reg_244][3  ( .D(D_3), .E(n6435), .C(wclk), .QN(n285) );
  DFE1 \mem_reg_244][2  ( .D(D_2), .E(n6435), .C(wclk), .QN(n286) );
  DFE1 \mem_reg_244][1  ( .D(D_1), .E(n6435), .C(wclk), .QN(n287) );
  DFE1 \mem_reg_244][0  ( .D(D_0), .E(n6435), .C(wclk), .QN(n288) );
  DFE1 \mem_reg_240][23  ( .D(D_23), .E(n6416), .C(wclk), .QN(n361) );
  DFE1 \mem_reg_240][22  ( .D(D_22), .E(n6416), .C(wclk), .QN(n362) );
  DFE1 \mem_reg_240][21  ( .D(D_21), .E(n6416), .C(wclk), .QN(n363) );
  DFE1 \mem_reg_240][20  ( .D(D_20), .E(n6416), .C(wclk), .QN(n364) );
  DFE1 \mem_reg_240][19  ( .D(D_19), .E(n6416), .C(wclk), .QN(n365) );
  DFE1 \mem_reg_240][18  ( .D(D_18), .E(n6416), .C(wclk), .QN(n366) );
  DFE1 \mem_reg_240][17  ( .D(D_17), .E(n6416), .C(wclk), .QN(n367) );
  DFE1 \mem_reg_240][16  ( .D(D_16), .E(n6416), .C(wclk), .QN(n368) );
  DFE1 \mem_reg_240][15  ( .D(D_15), .E(n6416), .C(wclk), .QN(n369) );
  DFE1 \mem_reg_240][14  ( .D(D_14), .E(n6416), .C(wclk), .QN(n370) );
  DFE1 \mem_reg_240][13  ( .D(D_13), .E(n6416), .C(wclk), .QN(n371) );
  DFE1 \mem_reg_240][12  ( .D(D_12), .E(n6416), .C(wclk), .QN(n372) );
  DFE1 \mem_reg_240][11  ( .D(D_11), .E(n6416), .C(wclk), .QN(n373) );
  DFE1 \mem_reg_240][10  ( .D(D_10), .E(n6416), .C(wclk), .QN(n374) );
  DFE1 \mem_reg_240][9  ( .D(D_9), .E(n6416), .C(wclk), .QN(n375) );
  DFE1 \mem_reg_240][8  ( .D(D_8), .E(n6416), .C(wclk), .QN(n376) );
  DFE1 \mem_reg_240][7  ( .D(D_7), .E(n6416), .C(wclk), .QN(n377) );
  DFE1 \mem_reg_240][6  ( .D(D_6), .E(n6416), .C(wclk), .QN(n378) );
  DFE1 \mem_reg_240][5  ( .D(D_5), .E(n6416), .C(wclk), .QN(n379) );
  DFE1 \mem_reg_240][4  ( .D(D_4), .E(n6416), .C(wclk), .QN(n380) );
  DFE1 \mem_reg_240][3  ( .D(D_3), .E(n6416), .C(wclk), .QN(n381) );
  DFE1 \mem_reg_240][2  ( .D(D_2), .E(n6416), .C(wclk), .QN(n382) );
  DFE1 \mem_reg_240][1  ( .D(D_1), .E(n6416), .C(wclk), .QN(n383) );
  DFE1 \mem_reg_240][0  ( .D(D_0), .E(n6416), .C(wclk), .QN(n384) );
  DFE1 \mem_reg_249][23  ( .D(D_23), .E(n6199), .C(wclk), .QN(n145) );
  DFE1 \mem_reg_249][22  ( .D(D_22), .E(n6199), .C(wclk), .QN(n146) );
  DFE1 \mem_reg_249][21  ( .D(D_21), .E(n6199), .C(wclk), .QN(n147) );
  DFE1 \mem_reg_249][20  ( .D(D_20), .E(n6199), .C(wclk), .QN(n148) );
  DFE1 \mem_reg_249][19  ( .D(D_19), .E(n6199), .C(wclk), .QN(n149) );
  DFE1 \mem_reg_249][18  ( .D(D_18), .E(n6199), .C(wclk), .QN(n150) );
  DFE1 \mem_reg_249][17  ( .D(D_17), .E(n6199), .C(wclk), .QN(n151) );
  DFE1 \mem_reg_249][16  ( .D(D_16), .E(n6199), .C(wclk), .QN(n152) );
  DFE1 \mem_reg_249][15  ( .D(D_15), .E(n6199), .C(wclk), .QN(n153) );
  DFE1 \mem_reg_249][14  ( .D(D_14), .E(n6199), .C(wclk), .QN(n154) );
  DFE1 \mem_reg_249][13  ( .D(D_13), .E(n6199), .C(wclk), .QN(n155) );
  DFE1 \mem_reg_249][12  ( .D(D_12), .E(n6199), .C(wclk), .QN(n156) );
  DFE1 \mem_reg_249][11  ( .D(D_11), .E(n6199), .C(wclk), .QN(n157) );
  DFE1 \mem_reg_249][10  ( .D(D_10), .E(n6199), .C(wclk), .QN(n158) );
  DFE1 \mem_reg_249][9  ( .D(D_9), .E(n6199), .C(wclk), .QN(n159) );
  DFE1 \mem_reg_249][8  ( .D(D_8), .E(n6199), .C(wclk), .QN(n160) );
  DFE1 \mem_reg_249][7  ( .D(D_7), .E(n6199), .C(wclk), .QN(n161) );
  DFE1 \mem_reg_249][6  ( .D(D_6), .E(n6199), .C(wclk), .QN(n162) );
  DFE1 \mem_reg_249][5  ( .D(D_5), .E(n6199), .C(wclk), .QN(n163) );
  DFE1 \mem_reg_249][4  ( .D(D_4), .E(n6199), .C(wclk), .QN(n164) );
  DFE1 \mem_reg_249][3  ( .D(D_3), .E(n6199), .C(wclk), .QN(n165) );
  DFE1 \mem_reg_249][2  ( .D(D_2), .E(n6199), .C(wclk), .QN(n166) );
  DFE1 \mem_reg_249][1  ( .D(D_1), .E(n6199), .C(wclk), .QN(n167) );
  DFE1 \mem_reg_249][0  ( .D(D_0), .E(n6199), .C(wclk), .QN(n168) );
  DFE1 \mem_reg_245][23  ( .D(D_23), .E(n6448), .C(wclk), .QN(n241) );
  DFE1 \mem_reg_245][22  ( .D(D_22), .E(n6448), .C(wclk), .QN(n242) );
  DFE1 \mem_reg_245][21  ( .D(D_21), .E(n6448), .C(wclk), .QN(n243) );
  DFE1 \mem_reg_245][20  ( .D(D_20), .E(n6448), .C(wclk), .QN(n244) );
  DFE1 \mem_reg_245][19  ( .D(D_19), .E(n6448), .C(wclk), .QN(n245) );
  DFE1 \mem_reg_245][18  ( .D(D_18), .E(n6448), .C(wclk), .QN(n246) );
  DFE1 \mem_reg_245][17  ( .D(D_17), .E(n6448), .C(wclk), .QN(n247) );
  DFE1 \mem_reg_245][16  ( .D(D_16), .E(n6448), .C(wclk), .QN(n248) );
  DFE1 \mem_reg_245][15  ( .D(D_15), .E(n6448), .C(wclk), .QN(n249) );
  DFE1 \mem_reg_245][14  ( .D(D_14), .E(n6448), .C(wclk), .QN(n250) );
  DFE1 \mem_reg_245][13  ( .D(D_13), .E(n6448), .C(wclk), .QN(n251) );
  DFE1 \mem_reg_245][12  ( .D(D_12), .E(n6448), .C(wclk), .QN(n252) );
  DFE1 \mem_reg_245][11  ( .D(D_11), .E(n6448), .C(wclk), .QN(n253) );
  DFE1 \mem_reg_245][10  ( .D(D_10), .E(n6448), .C(wclk), .QN(n254) );
  DFE1 \mem_reg_245][9  ( .D(D_9), .E(n6448), .C(wclk), .QN(n255) );
  DFE1 \mem_reg_245][8  ( .D(D_8), .E(n6448), .C(wclk), .QN(n256) );
  DFE1 \mem_reg_245][7  ( .D(D_7), .E(n6448), .C(wclk), .QN(n257) );
  DFE1 \mem_reg_245][6  ( .D(D_6), .E(n6448), .C(wclk), .QN(n258) );
  DFE1 \mem_reg_245][5  ( .D(D_5), .E(n6448), .C(wclk), .QN(n259) );
  DFE1 \mem_reg_245][4  ( .D(D_4), .E(n6448), .C(wclk), .QN(n260) );
  DFE1 \mem_reg_245][3  ( .D(D_3), .E(n6448), .C(wclk), .QN(n261) );
  DFE1 \mem_reg_245][2  ( .D(D_2), .E(n6448), .C(wclk), .QN(n262) );
  DFE1 \mem_reg_245][1  ( .D(D_1), .E(n6448), .C(wclk), .QN(n263) );
  DFE1 \mem_reg_245][0  ( .D(D_0), .E(n6448), .C(wclk), .QN(n264) );
  DFE1 \mem_reg_241][23  ( .D(D_23), .E(n6417), .C(wclk), .QN(n337) );
  DFE1 \mem_reg_241][22  ( .D(D_22), .E(n6417), .C(wclk), .QN(n338) );
  DFE1 \mem_reg_241][21  ( .D(D_21), .E(n6417), .C(wclk), .QN(n339) );
  DFE1 \mem_reg_241][20  ( .D(D_20), .E(n6417), .C(wclk), .QN(n340) );
  DFE1 \mem_reg_241][19  ( .D(D_19), .E(n6417), .C(wclk), .QN(n341) );
  DFE1 \mem_reg_241][18  ( .D(D_18), .E(n6417), .C(wclk), .QN(n342) );
  DFE1 \mem_reg_241][17  ( .D(D_17), .E(n6417), .C(wclk), .QN(n343) );
  DFE1 \mem_reg_241][16  ( .D(D_16), .E(n6417), .C(wclk), .QN(n344) );
  DFE1 \mem_reg_241][15  ( .D(D_15), .E(n6417), .C(wclk), .QN(n345) );
  DFE1 \mem_reg_241][14  ( .D(D_14), .E(n6417), .C(wclk), .QN(n346) );
  DFE1 \mem_reg_241][13  ( .D(D_13), .E(n6417), .C(wclk), .QN(n347) );
  DFE1 \mem_reg_241][12  ( .D(D_12), .E(n6417), .C(wclk), .QN(n348) );
  DFE1 \mem_reg_241][11  ( .D(D_11), .E(n6417), .C(wclk), .QN(n349) );
  DFE1 \mem_reg_241][10  ( .D(D_10), .E(n6417), .C(wclk), .QN(n350) );
  DFE1 \mem_reg_241][9  ( .D(D_9), .E(n6417), .C(wclk), .QN(n351) );
  DFE1 \mem_reg_241][8  ( .D(D_8), .E(n6417), .C(wclk), .QN(n352) );
  DFE1 \mem_reg_241][7  ( .D(D_7), .E(n6417), .C(wclk), .QN(n353) );
  DFE1 \mem_reg_241][6  ( .D(D_6), .E(n6417), .C(wclk), .QN(n354) );
  DFE1 \mem_reg_241][5  ( .D(D_5), .E(n6417), .C(wclk), .QN(n355) );
  DFE1 \mem_reg_241][4  ( .D(D_4), .E(n6417), .C(wclk), .QN(n356) );
  DFE1 \mem_reg_241][3  ( .D(D_3), .E(n6417), .C(wclk), .QN(n357) );
  DFE1 \mem_reg_241][2  ( .D(D_2), .E(n6417), .C(wclk), .QN(n358) );
  DFE1 \mem_reg_241][1  ( .D(D_1), .E(n6417), .C(wclk), .QN(n359) );
  DFE1 \mem_reg_241][0  ( .D(D_0), .E(n6417), .C(wclk), .QN(n360) );
  DFE1 \mem_reg_251][23  ( .D(D_23), .E(n6241), .C(wclk), .QN(n97) );
  DFE1 \mem_reg_251][22  ( .D(D_22), .E(n6241), .C(wclk), .QN(n98) );
  DFE1 \mem_reg_251][21  ( .D(D_21), .E(n6241), .C(wclk), .QN(n99) );
  DFE1 \mem_reg_251][20  ( .D(D_20), .E(n6241), .C(wclk), .QN(n100) );
  DFE1 \mem_reg_251][19  ( .D(D_19), .E(n6241), .C(wclk), .QN(n101) );
  DFE1 \mem_reg_251][18  ( .D(D_18), .E(n6241), .C(wclk), .QN(n102) );
  DFE1 \mem_reg_251][17  ( .D(D_17), .E(n6241), .C(wclk), .QN(n103) );
  DFE1 \mem_reg_251][16  ( .D(D_16), .E(n6241), .C(wclk), .QN(n104) );
  DFE1 \mem_reg_251][15  ( .D(D_15), .E(n6241), .C(wclk), .QN(n105) );
  DFE1 \mem_reg_251][14  ( .D(D_14), .E(n6241), .C(wclk), .QN(n106) );
  DFE1 \mem_reg_251][13  ( .D(D_13), .E(n6241), .C(wclk), .QN(n107) );
  DFE1 \mem_reg_251][12  ( .D(D_12), .E(n6241), .C(wclk), .QN(n108) );
  DFE1 \mem_reg_251][11  ( .D(D_11), .E(n6241), .C(wclk), .QN(n109) );
  DFE1 \mem_reg_251][10  ( .D(D_10), .E(n6241), .C(wclk), .QN(n110) );
  DFE1 \mem_reg_251][9  ( .D(D_9), .E(n6241), .C(wclk), .QN(n111) );
  DFE1 \mem_reg_251][8  ( .D(D_8), .E(n6241), .C(wclk), .QN(n112) );
  DFE1 \mem_reg_251][7  ( .D(D_7), .E(n6241), .C(wclk), .QN(n113) );
  DFE1 \mem_reg_251][6  ( .D(D_6), .E(n6241), .C(wclk), .QN(n114) );
  DFE1 \mem_reg_251][5  ( .D(D_5), .E(n6241), .C(wclk), .QN(n115) );
  DFE1 \mem_reg_251][4  ( .D(D_4), .E(n6241), .C(wclk), .QN(n116) );
  DFE1 \mem_reg_251][3  ( .D(D_3), .E(n6241), .C(wclk), .QN(n117) );
  DFE1 \mem_reg_251][2  ( .D(D_2), .E(n6241), .C(wclk), .QN(n118) );
  DFE1 \mem_reg_251][1  ( .D(D_1), .E(n6241), .C(wclk), .QN(n119) );
  DFE1 \mem_reg_251][0  ( .D(D_0), .E(n6241), .C(wclk), .QN(n120) );
  DFE1 \mem_reg_250][23  ( .D(D_23), .E(n6223), .C(wclk), .QN(n121) );
  DFE1 \mem_reg_250][22  ( .D(D_22), .E(n6223), .C(wclk), .QN(n122) );
  DFE1 \mem_reg_250][21  ( .D(D_21), .E(n6223), .C(wclk), .QN(n123) );
  DFE1 \mem_reg_250][20  ( .D(D_20), .E(n6223), .C(wclk), .QN(n124) );
  DFE1 \mem_reg_250][19  ( .D(D_19), .E(n6223), .C(wclk), .QN(n125) );
  DFE1 \mem_reg_250][18  ( .D(D_18), .E(n6223), .C(wclk), .QN(n126) );
  DFE1 \mem_reg_250][17  ( .D(D_17), .E(n6223), .C(wclk), .QN(n127) );
  DFE1 \mem_reg_250][16  ( .D(D_16), .E(n6223), .C(wclk), .QN(n128) );
  DFE1 \mem_reg_250][15  ( .D(D_15), .E(n6223), .C(wclk), .QN(n129) );
  DFE1 \mem_reg_250][14  ( .D(D_14), .E(n6223), .C(wclk), .QN(n130) );
  DFE1 \mem_reg_250][13  ( .D(D_13), .E(n6223), .C(wclk), .QN(n131) );
  DFE1 \mem_reg_250][12  ( .D(D_12), .E(n6223), .C(wclk), .QN(n132) );
  DFE1 \mem_reg_250][11  ( .D(D_11), .E(n6223), .C(wclk), .QN(n133) );
  DFE1 \mem_reg_250][10  ( .D(D_10), .E(n6223), .C(wclk), .QN(n134) );
  DFE1 \mem_reg_250][9  ( .D(D_9), .E(n6223), .C(wclk), .QN(n135) );
  DFE1 \mem_reg_250][8  ( .D(D_8), .E(n6223), .C(wclk), .QN(n136) );
  DFE1 \mem_reg_250][7  ( .D(D_7), .E(n6223), .C(wclk), .QN(n137) );
  DFE1 \mem_reg_250][6  ( .D(D_6), .E(n6223), .C(wclk), .QN(n138) );
  DFE1 \mem_reg_250][5  ( .D(D_5), .E(n6223), .C(wclk), .QN(n139) );
  DFE1 \mem_reg_250][4  ( .D(D_4), .E(n6223), .C(wclk), .QN(n140) );
  DFE1 \mem_reg_250][3  ( .D(D_3), .E(n6223), .C(wclk), .QN(n141) );
  DFE1 \mem_reg_250][2  ( .D(D_2), .E(n6223), .C(wclk), .QN(n142) );
  DFE1 \mem_reg_250][1  ( .D(D_1), .E(n6223), .C(wclk), .QN(n143) );
  DFE1 \mem_reg_250][0  ( .D(D_0), .E(n6223), .C(wclk), .QN(n144) );
  DFE1 \mem_reg_253][23  ( .D(D_23), .E(n6265), .C(wclk), .QN(n49) );
  DFE1 \mem_reg_253][22  ( .D(D_22), .E(n6265), .C(wclk), .QN(n50) );
  DFE1 \mem_reg_253][21  ( .D(D_21), .E(n6265), .C(wclk), .QN(n51) );
  DFE1 \mem_reg_253][20  ( .D(D_20), .E(n6265), .C(wclk), .QN(n52) );
  DFE1 \mem_reg_253][19  ( .D(D_19), .E(n6265), .C(wclk), .QN(n53) );
  DFE1 \mem_reg_253][18  ( .D(D_18), .E(n6265), .C(wclk), .QN(n54) );
  DFE1 \mem_reg_253][17  ( .D(D_17), .E(n6265), .C(wclk), .QN(n55) );
  DFE1 \mem_reg_253][16  ( .D(D_16), .E(n6265), .C(wclk), .QN(n56) );
  DFE1 \mem_reg_253][15  ( .D(D_15), .E(n6265), .C(wclk), .QN(n57) );
  DFE1 \mem_reg_253][14  ( .D(D_14), .E(n6265), .C(wclk), .QN(n58) );
  DFE1 \mem_reg_253][13  ( .D(D_13), .E(n6265), .C(wclk), .QN(n59) );
  DFE1 \mem_reg_253][12  ( .D(D_12), .E(n6265), .C(wclk), .QN(n60) );
  DFE1 \mem_reg_253][11  ( .D(D_11), .E(n6265), .C(wclk), .QN(n61) );
  DFE1 \mem_reg_253][10  ( .D(D_10), .E(n6265), .C(wclk), .QN(n62) );
  DFE1 \mem_reg_253][9  ( .D(D_9), .E(n6265), .C(wclk), .QN(n63) );
  DFE1 \mem_reg_253][8  ( .D(D_8), .E(n6265), .C(wclk), .QN(n64) );
  DFE1 \mem_reg_253][7  ( .D(D_7), .E(n6265), .C(wclk), .QN(n65) );
  DFE1 \mem_reg_253][6  ( .D(D_6), .E(n6265), .C(wclk), .QN(n66) );
  DFE1 \mem_reg_253][5  ( .D(D_5), .E(n6265), .C(wclk), .QN(n67) );
  DFE1 \mem_reg_253][4  ( .D(D_4), .E(n6265), .C(wclk), .QN(n68) );
  DFE1 \mem_reg_253][3  ( .D(D_3), .E(n6265), .C(wclk), .QN(n69) );
  DFE1 \mem_reg_253][2  ( .D(D_2), .E(n6265), .C(wclk), .QN(n70) );
  DFE1 \mem_reg_253][1  ( .D(D_1), .E(n6265), .C(wclk), .QN(n71) );
  DFE1 \mem_reg_253][0  ( .D(D_0), .E(n6265), .C(wclk), .QN(n72) );
  DFE1 \mem_reg_248][23  ( .D(D_23), .E(n6194), .C(wclk), .QN(n169) );
  DFE1 \mem_reg_248][22  ( .D(D_22), .E(n6194), .C(wclk), .QN(n170) );
  DFE1 \mem_reg_248][21  ( .D(D_21), .E(n6194), .C(wclk), .QN(n171) );
  DFE1 \mem_reg_248][20  ( .D(D_20), .E(n6194), .C(wclk), .QN(n172) );
  DFE1 \mem_reg_248][19  ( .D(D_19), .E(n6194), .C(wclk), .QN(n173) );
  DFE1 \mem_reg_248][18  ( .D(D_18), .E(n6194), .C(wclk), .QN(n174) );
  DFE1 \mem_reg_248][17  ( .D(D_17), .E(n6194), .C(wclk), .QN(n175) );
  DFE1 \mem_reg_248][16  ( .D(D_16), .E(n6194), .C(wclk), .QN(n176) );
  DFE1 \mem_reg_248][15  ( .D(D_15), .E(n6194), .C(wclk), .QN(n177) );
  DFE1 \mem_reg_248][14  ( .D(D_14), .E(n6194), .C(wclk), .QN(n178) );
  DFE1 \mem_reg_248][13  ( .D(D_13), .E(n6194), .C(wclk), .QN(n179) );
  DFE1 \mem_reg_248][12  ( .D(D_12), .E(n6194), .C(wclk), .QN(n180) );
  DFE1 \mem_reg_248][11  ( .D(D_11), .E(n6194), .C(wclk), .QN(n181) );
  DFE1 \mem_reg_248][10  ( .D(D_10), .E(n6194), .C(wclk), .QN(n182) );
  DFE1 \mem_reg_248][9  ( .D(D_9), .E(n6194), .C(wclk), .QN(n183) );
  DFE1 \mem_reg_248][8  ( .D(D_8), .E(n6194), .C(wclk), .QN(n184) );
  DFE1 \mem_reg_248][7  ( .D(D_7), .E(n6194), .C(wclk), .QN(n185) );
  DFE1 \mem_reg_248][6  ( .D(D_6), .E(n6194), .C(wclk), .QN(n186) );
  DFE1 \mem_reg_248][5  ( .D(D_5), .E(n6194), .C(wclk), .QN(n187) );
  DFE1 \mem_reg_248][4  ( .D(D_4), .E(n6194), .C(wclk), .QN(n188) );
  DFE1 \mem_reg_248][3  ( .D(D_3), .E(n6194), .C(wclk), .QN(n189) );
  DFE1 \mem_reg_248][2  ( .D(D_2), .E(n6194), .C(wclk), .QN(n190) );
  DFE1 \mem_reg_248][1  ( .D(D_1), .E(n6194), .C(wclk), .QN(n191) );
  DFE1 \mem_reg_248][0  ( .D(D_0), .E(n6194), .C(wclk), .QN(n192) );
  DFE1 \mem_reg_71][23  ( .D(D_23), .E(n6216), .C(wclk), .QN(n4417) );
  DFE1 \mem_reg_71][22  ( .D(D_22), .E(n6216), .C(wclk), .QN(n4418) );
  DFE1 \mem_reg_71][21  ( .D(D_21), .E(n6216), .C(wclk), .QN(n4419) );
  DFE1 \mem_reg_71][20  ( .D(D_20), .E(n6216), .C(wclk), .QN(n4420) );
  DFE1 \mem_reg_71][19  ( .D(D_19), .E(n6216), .C(wclk), .QN(n4421) );
  DFE1 \mem_reg_71][18  ( .D(D_18), .E(n6216), .C(wclk), .QN(n4422) );
  DFE1 \mem_reg_71][17  ( .D(D_17), .E(n6216), .C(wclk), .QN(n4423) );
  DFE1 \mem_reg_71][16  ( .D(D_16), .E(n6216), .C(wclk), .QN(n4424) );
  DFE1 \mem_reg_71][15  ( .D(D_15), .E(n6216), .C(wclk), .QN(n4425) );
  DFE1 \mem_reg_71][14  ( .D(D_14), .E(n6216), .C(wclk), .QN(n4426) );
  DFE1 \mem_reg_71][13  ( .D(D_13), .E(n6216), .C(wclk), .QN(n4427) );
  DFE1 \mem_reg_71][12  ( .D(D_12), .E(n6216), .C(wclk), .QN(n4428) );
  DFE1 \mem_reg_71][11  ( .D(D_11), .E(n6216), .C(wclk), .QN(n4429) );
  DFE1 \mem_reg_71][10  ( .D(D_10), .E(n6216), .C(wclk), .QN(n4430) );
  DFE1 \mem_reg_71][9  ( .D(D_9), .E(n6216), .C(wclk), .QN(n4431) );
  DFE1 \mem_reg_71][8  ( .D(D_8), .E(n6216), .C(wclk), .QN(n4432) );
  DFE1 \mem_reg_71][7  ( .D(D_7), .E(n6216), .C(wclk), .QN(n4433) );
  DFE1 \mem_reg_71][6  ( .D(D_6), .E(n6216), .C(wclk), .QN(n4434) );
  DFE1 \mem_reg_71][5  ( .D(D_5), .E(n6216), .C(wclk), .QN(n4435) );
  DFE1 \mem_reg_71][4  ( .D(D_4), .E(n6216), .C(wclk), .QN(n4436) );
  DFE1 \mem_reg_71][3  ( .D(D_3), .E(n6216), .C(wclk), .QN(n4437) );
  DFE1 \mem_reg_71][2  ( .D(D_2), .E(n6216), .C(wclk), .QN(n4438) );
  DFE1 \mem_reg_71][1  ( .D(D_1), .E(n6216), .C(wclk), .QN(n4439) );
  DFE1 \mem_reg_71][0  ( .D(D_0), .E(n6216), .C(wclk), .QN(n4440) );
  DFE1 \mem_reg_70][23  ( .D(D_23), .E(n6214), .C(wclk), .QN(n4441) );
  DFE1 \mem_reg_70][22  ( .D(D_22), .E(n6214), .C(wclk), .QN(n4442) );
  DFE1 \mem_reg_70][21  ( .D(D_21), .E(n6214), .C(wclk), .QN(n4443) );
  DFE1 \mem_reg_70][20  ( .D(D_20), .E(n6214), .C(wclk), .QN(n4444) );
  DFE1 \mem_reg_70][19  ( .D(D_19), .E(n6214), .C(wclk), .QN(n4445) );
  DFE1 \mem_reg_70][18  ( .D(D_18), .E(n6214), .C(wclk), .QN(n4446) );
  DFE1 \mem_reg_70][17  ( .D(D_17), .E(n6214), .C(wclk), .QN(n4447) );
  DFE1 \mem_reg_70][16  ( .D(D_16), .E(n6214), .C(wclk), .QN(n4448) );
  DFE1 \mem_reg_70][15  ( .D(D_15), .E(n6214), .C(wclk), .QN(n4449) );
  DFE1 \mem_reg_70][14  ( .D(D_14), .E(n6214), .C(wclk), .QN(n4450) );
  DFE1 \mem_reg_70][13  ( .D(D_13), .E(n6214), .C(wclk), .QN(n4451) );
  DFE1 \mem_reg_70][12  ( .D(D_12), .E(n6214), .C(wclk), .QN(n4452) );
  DFE1 \mem_reg_70][11  ( .D(D_11), .E(n6214), .C(wclk), .QN(n4453) );
  DFE1 \mem_reg_70][10  ( .D(D_10), .E(n6214), .C(wclk), .QN(n4454) );
  DFE1 \mem_reg_70][9  ( .D(D_9), .E(n6214), .C(wclk), .QN(n4455) );
  DFE1 \mem_reg_70][8  ( .D(D_8), .E(n6214), .C(wclk), .QN(n4456) );
  DFE1 \mem_reg_70][7  ( .D(D_7), .E(n6214), .C(wclk), .QN(n4457) );
  DFE1 \mem_reg_70][6  ( .D(D_6), .E(n6214), .C(wclk), .QN(n4458) );
  DFE1 \mem_reg_70][5  ( .D(D_5), .E(n6214), .C(wclk), .QN(n4459) );
  DFE1 \mem_reg_70][4  ( .D(D_4), .E(n6214), .C(wclk), .QN(n4460) );
  DFE1 \mem_reg_70][3  ( .D(D_3), .E(n6214), .C(wclk), .QN(n4461) );
  DFE1 \mem_reg_70][2  ( .D(D_2), .E(n6214), .C(wclk), .QN(n4462) );
  DFE1 \mem_reg_70][1  ( .D(D_1), .E(n6214), .C(wclk), .QN(n4463) );
  DFE1 \mem_reg_70][0  ( .D(D_0), .E(n6214), .C(wclk), .QN(n4464) );
  DFE1 \mem_reg_67][23  ( .D(D_23), .E(n6208), .C(wclk), .QN(n4513) );
  DFE1 \mem_reg_67][22  ( .D(D_22), .E(n6208), .C(wclk), .QN(n4514) );
  DFE1 \mem_reg_67][21  ( .D(D_21), .E(n6208), .C(wclk), .QN(n4515) );
  DFE1 \mem_reg_67][20  ( .D(D_20), .E(n6208), .C(wclk), .QN(n4516) );
  DFE1 \mem_reg_67][19  ( .D(D_19), .E(n6208), .C(wclk), .QN(n4517) );
  DFE1 \mem_reg_67][18  ( .D(D_18), .E(n6208), .C(wclk), .QN(n4518) );
  DFE1 \mem_reg_67][17  ( .D(D_17), .E(n6208), .C(wclk), .QN(n4519) );
  DFE1 \mem_reg_67][16  ( .D(D_16), .E(n6208), .C(wclk), .QN(n4520) );
  DFE1 \mem_reg_67][15  ( .D(D_15), .E(n6208), .C(wclk), .QN(n4521) );
  DFE1 \mem_reg_67][14  ( .D(D_14), .E(n6208), .C(wclk), .QN(n4522) );
  DFE1 \mem_reg_67][13  ( .D(D_13), .E(n6208), .C(wclk), .QN(n4523) );
  DFE1 \mem_reg_67][12  ( .D(D_12), .E(n6208), .C(wclk), .QN(n4524) );
  DFE1 \mem_reg_67][11  ( .D(D_11), .E(n6208), .C(wclk), .QN(n4525) );
  DFE1 \mem_reg_67][10  ( .D(D_10), .E(n6208), .C(wclk), .QN(n4526) );
  DFE1 \mem_reg_67][9  ( .D(D_9), .E(n6208), .C(wclk), .QN(n4527) );
  DFE1 \mem_reg_67][8  ( .D(D_8), .E(n6208), .C(wclk), .QN(n4528) );
  DFE1 \mem_reg_67][7  ( .D(D_7), .E(n6208), .C(wclk), .QN(n4529) );
  DFE1 \mem_reg_67][6  ( .D(D_6), .E(n6208), .C(wclk), .QN(n4530) );
  DFE1 \mem_reg_67][5  ( .D(D_5), .E(n6208), .C(wclk), .QN(n4531) );
  DFE1 \mem_reg_67][4  ( .D(D_4), .E(n6208), .C(wclk), .QN(n4532) );
  DFE1 \mem_reg_67][3  ( .D(D_3), .E(n6208), .C(wclk), .QN(n4533) );
  DFE1 \mem_reg_67][2  ( .D(D_2), .E(n6208), .C(wclk), .QN(n4534) );
  DFE1 \mem_reg_67][1  ( .D(D_1), .E(n6208), .C(wclk), .QN(n4535) );
  DFE1 \mem_reg_67][0  ( .D(D_0), .E(n6208), .C(wclk), .QN(n4536) );
  DFE1 \mem_reg_66][23  ( .D(D_23), .E(n6206), .C(wclk), .QN(n4537) );
  DFE1 \mem_reg_66][22  ( .D(D_22), .E(n6206), .C(wclk), .QN(n4538) );
  DFE1 \mem_reg_66][21  ( .D(D_21), .E(n6206), .C(wclk), .QN(n4539) );
  DFE1 \mem_reg_66][20  ( .D(D_20), .E(n6206), .C(wclk), .QN(n4540) );
  DFE1 \mem_reg_66][19  ( .D(D_19), .E(n6206), .C(wclk), .QN(n4541) );
  DFE1 \mem_reg_66][18  ( .D(D_18), .E(n6206), .C(wclk), .QN(n4542) );
  DFE1 \mem_reg_66][17  ( .D(D_17), .E(n6206), .C(wclk), .QN(n4543) );
  DFE1 \mem_reg_66][16  ( .D(D_16), .E(n6206), .C(wclk), .QN(n4544) );
  DFE1 \mem_reg_66][15  ( .D(D_15), .E(n6206), .C(wclk), .QN(n4545) );
  DFE1 \mem_reg_66][14  ( .D(D_14), .E(n6206), .C(wclk), .QN(n4546) );
  DFE1 \mem_reg_66][13  ( .D(D_13), .E(n6206), .C(wclk), .QN(n4547) );
  DFE1 \mem_reg_66][12  ( .D(D_12), .E(n6206), .C(wclk), .QN(n4548) );
  DFE1 \mem_reg_66][11  ( .D(D_11), .E(n6206), .C(wclk), .QN(n4549) );
  DFE1 \mem_reg_66][10  ( .D(D_10), .E(n6206), .C(wclk), .QN(n4550) );
  DFE1 \mem_reg_66][9  ( .D(D_9), .E(n6206), .C(wclk), .QN(n4551) );
  DFE1 \mem_reg_66][8  ( .D(D_8), .E(n6206), .C(wclk), .QN(n4552) );
  DFE1 \mem_reg_66][7  ( .D(D_7), .E(n6206), .C(wclk), .QN(n4553) );
  DFE1 \mem_reg_66][6  ( .D(D_6), .E(n6206), .C(wclk), .QN(n4554) );
  DFE1 \mem_reg_66][5  ( .D(D_5), .E(n6206), .C(wclk), .QN(n4555) );
  DFE1 \mem_reg_66][4  ( .D(D_4), .E(n6206), .C(wclk), .QN(n4556) );
  DFE1 \mem_reg_66][3  ( .D(D_3), .E(n6206), .C(wclk), .QN(n4557) );
  DFE1 \mem_reg_66][2  ( .D(D_2), .E(n6206), .C(wclk), .QN(n4558) );
  DFE1 \mem_reg_66][1  ( .D(D_1), .E(n6206), .C(wclk), .QN(n4559) );
  DFE1 \mem_reg_66][0  ( .D(D_0), .E(n6206), .C(wclk), .QN(n4560) );
  DFE1 \mem_reg_76][23  ( .D(D_23), .E(n6228), .C(wclk), .QN(n4297) );
  DFE1 \mem_reg_76][22  ( .D(D_22), .E(n6228), .C(wclk), .QN(n4298) );
  DFE1 \mem_reg_76][21  ( .D(D_21), .E(n6228), .C(wclk), .QN(n4299) );
  DFE1 \mem_reg_76][20  ( .D(D_20), .E(n6228), .C(wclk), .QN(n4300) );
  DFE1 \mem_reg_76][19  ( .D(D_19), .E(n6228), .C(wclk), .QN(n4301) );
  DFE1 \mem_reg_76][18  ( .D(D_18), .E(n6228), .C(wclk), .QN(n4302) );
  DFE1 \mem_reg_76][17  ( .D(D_17), .E(n6228), .C(wclk), .QN(n4303) );
  DFE1 \mem_reg_76][16  ( .D(D_16), .E(n6228), .C(wclk), .QN(n4304) );
  DFE1 \mem_reg_76][15  ( .D(D_15), .E(n6228), .C(wclk), .QN(n4305) );
  DFE1 \mem_reg_76][14  ( .D(D_14), .E(n6228), .C(wclk), .QN(n4306) );
  DFE1 \mem_reg_76][13  ( .D(D_13), .E(n6228), .C(wclk), .QN(n4307) );
  DFE1 \mem_reg_76][12  ( .D(D_12), .E(n6228), .C(wclk), .QN(n4308) );
  DFE1 \mem_reg_76][11  ( .D(D_11), .E(n6228), .C(wclk), .QN(n4309) );
  DFE1 \mem_reg_76][10  ( .D(D_10), .E(n6228), .C(wclk), .QN(n4310) );
  DFE1 \mem_reg_76][9  ( .D(D_9), .E(n6228), .C(wclk), .QN(n4311) );
  DFE1 \mem_reg_76][8  ( .D(D_8), .E(n6228), .C(wclk), .QN(n4312) );
  DFE1 \mem_reg_76][7  ( .D(D_7), .E(n6228), .C(wclk), .QN(n4313) );
  DFE1 \mem_reg_76][6  ( .D(D_6), .E(n6228), .C(wclk), .QN(n4314) );
  DFE1 \mem_reg_76][5  ( .D(D_5), .E(n6228), .C(wclk), .QN(n4315) );
  DFE1 \mem_reg_76][4  ( .D(D_4), .E(n6228), .C(wclk), .QN(n4316) );
  DFE1 \mem_reg_76][3  ( .D(D_3), .E(n6228), .C(wclk), .QN(n4317) );
  DFE1 \mem_reg_76][2  ( .D(D_2), .E(n6228), .C(wclk), .QN(n4318) );
  DFE1 \mem_reg_76][1  ( .D(D_1), .E(n6228), .C(wclk), .QN(n4319) );
  DFE1 \mem_reg_76][0  ( .D(D_0), .E(n6228), .C(wclk), .QN(n4320) );
  DFE1 \mem_reg_68][23  ( .D(D_23), .E(n6210), .C(wclk), .QN(n4489) );
  DFE1 \mem_reg_68][22  ( .D(D_22), .E(n6210), .C(wclk), .QN(n4490) );
  DFE1 \mem_reg_68][21  ( .D(D_21), .E(n6210), .C(wclk), .QN(n4491) );
  DFE1 \mem_reg_68][20  ( .D(D_20), .E(n6210), .C(wclk), .QN(n4492) );
  DFE1 \mem_reg_68][19  ( .D(D_19), .E(n6210), .C(wclk), .QN(n4493) );
  DFE1 \mem_reg_68][18  ( .D(D_18), .E(n6210), .C(wclk), .QN(n4494) );
  DFE1 \mem_reg_68][17  ( .D(D_17), .E(n6210), .C(wclk), .QN(n4495) );
  DFE1 \mem_reg_68][16  ( .D(D_16), .E(n6210), .C(wclk), .QN(n4496) );
  DFE1 \mem_reg_68][15  ( .D(D_15), .E(n6210), .C(wclk), .QN(n4497) );
  DFE1 \mem_reg_68][14  ( .D(D_14), .E(n6210), .C(wclk), .QN(n4498) );
  DFE1 \mem_reg_68][13  ( .D(D_13), .E(n6210), .C(wclk), .QN(n4499) );
  DFE1 \mem_reg_68][12  ( .D(D_12), .E(n6210), .C(wclk), .QN(n4500) );
  DFE1 \mem_reg_68][11  ( .D(D_11), .E(n6210), .C(wclk), .QN(n4501) );
  DFE1 \mem_reg_68][10  ( .D(D_10), .E(n6210), .C(wclk), .QN(n4502) );
  DFE1 \mem_reg_68][9  ( .D(D_9), .E(n6210), .C(wclk), .QN(n4503) );
  DFE1 \mem_reg_68][8  ( .D(D_8), .E(n6210), .C(wclk), .QN(n4504) );
  DFE1 \mem_reg_68][7  ( .D(D_7), .E(n6210), .C(wclk), .QN(n4505) );
  DFE1 \mem_reg_68][6  ( .D(D_6), .E(n6210), .C(wclk), .QN(n4506) );
  DFE1 \mem_reg_68][5  ( .D(D_5), .E(n6210), .C(wclk), .QN(n4507) );
  DFE1 \mem_reg_68][4  ( .D(D_4), .E(n6210), .C(wclk), .QN(n4508) );
  DFE1 \mem_reg_68][3  ( .D(D_3), .E(n6210), .C(wclk), .QN(n4509) );
  DFE1 \mem_reg_68][2  ( .D(D_2), .E(n6210), .C(wclk), .QN(n4510) );
  DFE1 \mem_reg_68][1  ( .D(D_1), .E(n6210), .C(wclk), .QN(n4511) );
  DFE1 \mem_reg_68][0  ( .D(D_0), .E(n6210), .C(wclk), .QN(n4512) );
  DFE1 \mem_reg_69][23  ( .D(D_23), .E(n6212), .C(wclk), .QN(n4465) );
  DFE1 \mem_reg_69][22  ( .D(D_22), .E(n6212), .C(wclk), .QN(n4466) );
  DFE1 \mem_reg_69][21  ( .D(D_21), .E(n6212), .C(wclk), .QN(n4467) );
  DFE1 \mem_reg_69][20  ( .D(D_20), .E(n6212), .C(wclk), .QN(n4468) );
  DFE1 \mem_reg_69][19  ( .D(D_19), .E(n6212), .C(wclk), .QN(n4469) );
  DFE1 \mem_reg_69][18  ( .D(D_18), .E(n6212), .C(wclk), .QN(n4470) );
  DFE1 \mem_reg_69][17  ( .D(D_17), .E(n6212), .C(wclk), .QN(n4471) );
  DFE1 \mem_reg_69][16  ( .D(D_16), .E(n6212), .C(wclk), .QN(n4472) );
  DFE1 \mem_reg_69][15  ( .D(D_15), .E(n6212), .C(wclk), .QN(n4473) );
  DFE1 \mem_reg_69][14  ( .D(D_14), .E(n6212), .C(wclk), .QN(n4474) );
  DFE1 \mem_reg_69][13  ( .D(D_13), .E(n6212), .C(wclk), .QN(n4475) );
  DFE1 \mem_reg_69][12  ( .D(D_12), .E(n6212), .C(wclk), .QN(n4476) );
  DFE1 \mem_reg_69][11  ( .D(D_11), .E(n6212), .C(wclk), .QN(n4477) );
  DFE1 \mem_reg_69][10  ( .D(D_10), .E(n6212), .C(wclk), .QN(n4478) );
  DFE1 \mem_reg_69][9  ( .D(D_9), .E(n6212), .C(wclk), .QN(n4479) );
  DFE1 \mem_reg_69][8  ( .D(D_8), .E(n6212), .C(wclk), .QN(n4480) );
  DFE1 \mem_reg_69][7  ( .D(D_7), .E(n6212), .C(wclk), .QN(n4481) );
  DFE1 \mem_reg_69][6  ( .D(D_6), .E(n6212), .C(wclk), .QN(n4482) );
  DFE1 \mem_reg_69][5  ( .D(D_5), .E(n6212), .C(wclk), .QN(n4483) );
  DFE1 \mem_reg_69][4  ( .D(D_4), .E(n6212), .C(wclk), .QN(n4484) );
  DFE1 \mem_reg_69][3  ( .D(D_3), .E(n6212), .C(wclk), .QN(n4485) );
  DFE1 \mem_reg_69][2  ( .D(D_2), .E(n6212), .C(wclk), .QN(n4486) );
  DFE1 \mem_reg_69][1  ( .D(D_1), .E(n6212), .C(wclk), .QN(n4487) );
  DFE1 \mem_reg_69][0  ( .D(D_0), .E(n6212), .C(wclk), .QN(n4488) );
  DFE1 \mem_reg_65][23  ( .D(D_23), .E(n6204), .C(wclk), .QN(n4561) );
  DFE1 \mem_reg_65][22  ( .D(D_22), .E(n6204), .C(wclk), .QN(n4562) );
  DFE1 \mem_reg_65][21  ( .D(D_21), .E(n6204), .C(wclk), .QN(n4563) );
  DFE1 \mem_reg_65][20  ( .D(D_20), .E(n6204), .C(wclk), .QN(n4564) );
  DFE1 \mem_reg_65][19  ( .D(D_19), .E(n6204), .C(wclk), .QN(n4565) );
  DFE1 \mem_reg_65][18  ( .D(D_18), .E(n6204), .C(wclk), .QN(n4566) );
  DFE1 \mem_reg_65][17  ( .D(D_17), .E(n6204), .C(wclk), .QN(n4567) );
  DFE1 \mem_reg_65][16  ( .D(D_16), .E(n6204), .C(wclk), .QN(n4568) );
  DFE1 \mem_reg_65][15  ( .D(D_15), .E(n6204), .C(wclk), .QN(n4569) );
  DFE1 \mem_reg_65][14  ( .D(D_14), .E(n6204), .C(wclk), .QN(n4570) );
  DFE1 \mem_reg_65][13  ( .D(D_13), .E(n6204), .C(wclk), .QN(n4571) );
  DFE1 \mem_reg_65][12  ( .D(D_12), .E(n6204), .C(wclk), .QN(n4572) );
  DFE1 \mem_reg_65][11  ( .D(D_11), .E(n6204), .C(wclk), .QN(n4573) );
  DFE1 \mem_reg_65][10  ( .D(D_10), .E(n6204), .C(wclk), .QN(n4574) );
  DFE1 \mem_reg_65][9  ( .D(D_9), .E(n6204), .C(wclk), .QN(n4575) );
  DFE1 \mem_reg_65][8  ( .D(D_8), .E(n6204), .C(wclk), .QN(n4576) );
  DFE1 \mem_reg_65][7  ( .D(D_7), .E(n6204), .C(wclk), .QN(n4577) );
  DFE1 \mem_reg_65][6  ( .D(D_6), .E(n6204), .C(wclk), .QN(n4578) );
  DFE1 \mem_reg_65][5  ( .D(D_5), .E(n6204), .C(wclk), .QN(n4579) );
  DFE1 \mem_reg_65][4  ( .D(D_4), .E(n6204), .C(wclk), .QN(n4580) );
  DFE1 \mem_reg_65][3  ( .D(D_3), .E(n6204), .C(wclk), .QN(n4581) );
  DFE1 \mem_reg_65][2  ( .D(D_2), .E(n6204), .C(wclk), .QN(n4582) );
  DFE1 \mem_reg_65][1  ( .D(D_1), .E(n6204), .C(wclk), .QN(n4583) );
  DFE1 \mem_reg_65][0  ( .D(D_0), .E(n6204), .C(wclk), .QN(n4584) );
  DFE1 \mem_reg_75][23  ( .D(D_23), .E(n6226), .C(wclk), .QN(n4321) );
  DFE1 \mem_reg_75][22  ( .D(D_22), .E(n6226), .C(wclk), .QN(n4322) );
  DFE1 \mem_reg_75][21  ( .D(D_21), .E(n6226), .C(wclk), .QN(n4323) );
  DFE1 \mem_reg_75][20  ( .D(D_20), .E(n6226), .C(wclk), .QN(n4324) );
  DFE1 \mem_reg_75][19  ( .D(D_19), .E(n6226), .C(wclk), .QN(n4325) );
  DFE1 \mem_reg_75][18  ( .D(D_18), .E(n6226), .C(wclk), .QN(n4326) );
  DFE1 \mem_reg_75][17  ( .D(D_17), .E(n6226), .C(wclk), .QN(n4327) );
  DFE1 \mem_reg_75][16  ( .D(D_16), .E(n6226), .C(wclk), .QN(n4328) );
  DFE1 \mem_reg_75][15  ( .D(D_15), .E(n6226), .C(wclk), .QN(n4329) );
  DFE1 \mem_reg_75][14  ( .D(D_14), .E(n6226), .C(wclk), .QN(n4330) );
  DFE1 \mem_reg_75][13  ( .D(D_13), .E(n6226), .C(wclk), .QN(n4331) );
  DFE1 \mem_reg_75][12  ( .D(D_12), .E(n6226), .C(wclk), .QN(n4332) );
  DFE1 \mem_reg_75][11  ( .D(D_11), .E(n6226), .C(wclk), .QN(n4333) );
  DFE1 \mem_reg_75][10  ( .D(D_10), .E(n6226), .C(wclk), .QN(n4334) );
  DFE1 \mem_reg_75][9  ( .D(D_9), .E(n6226), .C(wclk), .QN(n4335) );
  DFE1 \mem_reg_75][8  ( .D(D_8), .E(n6226), .C(wclk), .QN(n4336) );
  DFE1 \mem_reg_75][7  ( .D(D_7), .E(n6226), .C(wclk), .QN(n4337) );
  DFE1 \mem_reg_75][6  ( .D(D_6), .E(n6226), .C(wclk), .QN(n4338) );
  DFE1 \mem_reg_75][5  ( .D(D_5), .E(n6226), .C(wclk), .QN(n4339) );
  DFE1 \mem_reg_75][4  ( .D(D_4), .E(n6226), .C(wclk), .QN(n4340) );
  DFE1 \mem_reg_75][3  ( .D(D_3), .E(n6226), .C(wclk), .QN(n4341) );
  DFE1 \mem_reg_75][2  ( .D(D_2), .E(n6226), .C(wclk), .QN(n4342) );
  DFE1 \mem_reg_75][1  ( .D(D_1), .E(n6226), .C(wclk), .QN(n4343) );
  DFE1 \mem_reg_75][0  ( .D(D_0), .E(n6226), .C(wclk), .QN(n4344) );
  DFE1 \mem_reg_74][23  ( .D(D_23), .E(n6224), .C(wclk), .QN(n4345) );
  DFE1 \mem_reg_74][22  ( .D(D_22), .E(n6224), .C(wclk), .QN(n4346) );
  DFE1 \mem_reg_74][21  ( .D(D_21), .E(n6224), .C(wclk), .QN(n4347) );
  DFE1 \mem_reg_74][20  ( .D(D_20), .E(n6224), .C(wclk), .QN(n4348) );
  DFE1 \mem_reg_74][19  ( .D(D_19), .E(n6224), .C(wclk), .QN(n4349) );
  DFE1 \mem_reg_74][18  ( .D(D_18), .E(n6224), .C(wclk), .QN(n4350) );
  DFE1 \mem_reg_74][17  ( .D(D_17), .E(n6224), .C(wclk), .QN(n4351) );
  DFE1 \mem_reg_74][16  ( .D(D_16), .E(n6224), .C(wclk), .QN(n4352) );
  DFE1 \mem_reg_74][15  ( .D(D_15), .E(n6224), .C(wclk), .QN(n4353) );
  DFE1 \mem_reg_74][14  ( .D(D_14), .E(n6224), .C(wclk), .QN(n4354) );
  DFE1 \mem_reg_74][13  ( .D(D_13), .E(n6224), .C(wclk), .QN(n4355) );
  DFE1 \mem_reg_74][12  ( .D(D_12), .E(n6224), .C(wclk), .QN(n4356) );
  DFE1 \mem_reg_74][11  ( .D(D_11), .E(n6224), .C(wclk), .QN(n4357) );
  DFE1 \mem_reg_74][10  ( .D(D_10), .E(n6224), .C(wclk), .QN(n4358) );
  DFE1 \mem_reg_74][9  ( .D(D_9), .E(n6224), .C(wclk), .QN(n4359) );
  DFE1 \mem_reg_74][8  ( .D(D_8), .E(n6224), .C(wclk), .QN(n4360) );
  DFE1 \mem_reg_74][7  ( .D(D_7), .E(n6224), .C(wclk), .QN(n4361) );
  DFE1 \mem_reg_74][6  ( .D(D_6), .E(n6224), .C(wclk), .QN(n4362) );
  DFE1 \mem_reg_74][5  ( .D(D_5), .E(n6224), .C(wclk), .QN(n4363) );
  DFE1 \mem_reg_74][4  ( .D(D_4), .E(n6224), .C(wclk), .QN(n4364) );
  DFE1 \mem_reg_74][3  ( .D(D_3), .E(n6224), .C(wclk), .QN(n4365) );
  DFE1 \mem_reg_74][2  ( .D(D_2), .E(n6224), .C(wclk), .QN(n4366) );
  DFE1 \mem_reg_74][1  ( .D(D_1), .E(n6224), .C(wclk), .QN(n4367) );
  DFE1 \mem_reg_74][0  ( .D(D_0), .E(n6224), .C(wclk), .QN(n4368) );
  DFE1 \mem_reg_191][23  ( .D(D_23), .E(n6363), .C(wclk), .QN(n1537) );
  DFE1 \mem_reg_191][22  ( .D(D_22), .E(n6363), .C(wclk), .QN(n1538) );
  DFE1 \mem_reg_191][21  ( .D(D_21), .E(n6363), .C(wclk), .QN(n1539) );
  DFE1 \mem_reg_191][20  ( .D(D_20), .E(n6363), .C(wclk), .QN(n1540) );
  DFE1 \mem_reg_191][19  ( .D(D_19), .E(n6363), .C(wclk), .QN(n1541) );
  DFE1 \mem_reg_191][18  ( .D(D_18), .E(n6363), .C(wclk), .QN(n1542) );
  DFE1 \mem_reg_191][17  ( .D(D_17), .E(n6363), .C(wclk), .QN(n1543) );
  DFE1 \mem_reg_191][16  ( .D(D_16), .E(n6363), .C(wclk), .QN(n1544) );
  DFE1 \mem_reg_191][15  ( .D(D_15), .E(n6363), .C(wclk), .QN(n1545) );
  DFE1 \mem_reg_191][14  ( .D(D_14), .E(n6363), .C(wclk), .QN(n1546) );
  DFE1 \mem_reg_191][13  ( .D(D_13), .E(n6363), .C(wclk), .QN(n1547) );
  DFE1 \mem_reg_191][12  ( .D(D_12), .E(n6363), .C(wclk), .QN(n1548) );
  DFE1 \mem_reg_191][11  ( .D(D_11), .E(n6363), .C(wclk), .QN(n1549) );
  DFE1 \mem_reg_191][10  ( .D(D_10), .E(n6363), .C(wclk), .QN(n1550) );
  DFE1 \mem_reg_191][9  ( .D(D_9), .E(n6363), .C(wclk), .QN(n1551) );
  DFE1 \mem_reg_191][8  ( .D(D_8), .E(n6363), .C(wclk), .QN(n1552) );
  DFE1 \mem_reg_191][7  ( .D(D_7), .E(n6363), .C(wclk), .QN(n1553) );
  DFE1 \mem_reg_191][6  ( .D(D_6), .E(n6363), .C(wclk), .QN(n1554) );
  DFE1 \mem_reg_191][5  ( .D(D_5), .E(n6363), .C(wclk), .QN(n1555) );
  DFE1 \mem_reg_191][4  ( .D(D_4), .E(n6363), .C(wclk), .QN(n1556) );
  DFE1 \mem_reg_191][3  ( .D(D_3), .E(n6363), .C(wclk), .QN(n1557) );
  DFE1 \mem_reg_191][2  ( .D(D_2), .E(n6363), .C(wclk), .QN(n1558) );
  DFE1 \mem_reg_191][1  ( .D(D_1), .E(n6363), .C(wclk), .QN(n1559) );
  DFE1 \mem_reg_191][0  ( .D(D_0), .E(n6363), .C(wclk), .QN(n1560) );
  DFE1 \mem_reg_190][23  ( .D(D_23), .E(n6362), .C(wclk), .QN(n1561) );
  DFE1 \mem_reg_190][22  ( .D(D_22), .E(n6362), .C(wclk), .QN(n1562) );
  DFE1 \mem_reg_190][21  ( .D(D_21), .E(n6362), .C(wclk), .QN(n1563) );
  DFE1 \mem_reg_190][20  ( .D(D_20), .E(n6362), .C(wclk), .QN(n1564) );
  DFE1 \mem_reg_190][19  ( .D(D_19), .E(n6362), .C(wclk), .QN(n1565) );
  DFE1 \mem_reg_190][18  ( .D(D_18), .E(n6362), .C(wclk), .QN(n1566) );
  DFE1 \mem_reg_190][17  ( .D(D_17), .E(n6362), .C(wclk), .QN(n1567) );
  DFE1 \mem_reg_190][16  ( .D(D_16), .E(n6362), .C(wclk), .QN(n1568) );
  DFE1 \mem_reg_190][15  ( .D(D_15), .E(n6362), .C(wclk), .QN(n1569) );
  DFE1 \mem_reg_190][14  ( .D(D_14), .E(n6362), .C(wclk), .QN(n1570) );
  DFE1 \mem_reg_190][13  ( .D(D_13), .E(n6362), .C(wclk), .QN(n1571) );
  DFE1 \mem_reg_190][12  ( .D(D_12), .E(n6362), .C(wclk), .QN(n1572) );
  DFE1 \mem_reg_190][11  ( .D(D_11), .E(n6362), .C(wclk), .QN(n1573) );
  DFE1 \mem_reg_190][10  ( .D(D_10), .E(n6362), .C(wclk), .QN(n1574) );
  DFE1 \mem_reg_190][9  ( .D(D_9), .E(n6362), .C(wclk), .QN(n1575) );
  DFE1 \mem_reg_190][8  ( .D(D_8), .E(n6362), .C(wclk), .QN(n1576) );
  DFE1 \mem_reg_190][7  ( .D(D_7), .E(n6362), .C(wclk), .QN(n1577) );
  DFE1 \mem_reg_190][6  ( .D(D_6), .E(n6362), .C(wclk), .QN(n1578) );
  DFE1 \mem_reg_190][5  ( .D(D_5), .E(n6362), .C(wclk), .QN(n1579) );
  DFE1 \mem_reg_190][4  ( .D(D_4), .E(n6362), .C(wclk), .QN(n1580) );
  DFE1 \mem_reg_190][3  ( .D(D_3), .E(n6362), .C(wclk), .QN(n1581) );
  DFE1 \mem_reg_190][2  ( .D(D_2), .E(n6362), .C(wclk), .QN(n1582) );
  DFE1 \mem_reg_190][1  ( .D(D_1), .E(n6362), .C(wclk), .QN(n1583) );
  DFE1 \mem_reg_190][0  ( .D(D_0), .E(n6362), .C(wclk), .QN(n1584) );
  DFE1 \mem_reg_189][23  ( .D(D_23), .E(n6361), .C(wclk), .QN(n1585) );
  DFE1 \mem_reg_189][22  ( .D(D_22), .E(n6361), .C(wclk), .QN(n1586) );
  DFE1 \mem_reg_189][21  ( .D(D_21), .E(n6361), .C(wclk), .QN(n1587) );
  DFE1 \mem_reg_189][20  ( .D(D_20), .E(n6361), .C(wclk), .QN(n1588) );
  DFE1 \mem_reg_189][19  ( .D(D_19), .E(n6361), .C(wclk), .QN(n1589) );
  DFE1 \mem_reg_189][18  ( .D(D_18), .E(n6361), .C(wclk), .QN(n1590) );
  DFE1 \mem_reg_189][17  ( .D(D_17), .E(n6361), .C(wclk), .QN(n1591) );
  DFE1 \mem_reg_189][16  ( .D(D_16), .E(n6361), .C(wclk), .QN(n1592) );
  DFE1 \mem_reg_189][15  ( .D(D_15), .E(n6361), .C(wclk), .QN(n1593) );
  DFE1 \mem_reg_189][14  ( .D(D_14), .E(n6361), .C(wclk), .QN(n1594) );
  DFE1 \mem_reg_189][13  ( .D(D_13), .E(n6361), .C(wclk), .QN(n1595) );
  DFE1 \mem_reg_189][12  ( .D(D_12), .E(n6361), .C(wclk), .QN(n1596) );
  DFE1 \mem_reg_189][11  ( .D(D_11), .E(n6361), .C(wclk), .QN(n1597) );
  DFE1 \mem_reg_189][10  ( .D(D_10), .E(n6361), .C(wclk), .QN(n1598) );
  DFE1 \mem_reg_189][9  ( .D(D_9), .E(n6361), .C(wclk), .QN(n1599) );
  DFE1 \mem_reg_189][8  ( .D(D_8), .E(n6361), .C(wclk), .QN(n1600) );
  DFE1 \mem_reg_189][7  ( .D(D_7), .E(n6361), .C(wclk), .QN(n1601) );
  DFE1 \mem_reg_189][6  ( .D(D_6), .E(n6361), .C(wclk), .QN(n1602) );
  DFE1 \mem_reg_189][5  ( .D(D_5), .E(n6361), .C(wclk), .QN(n1603) );
  DFE1 \mem_reg_189][4  ( .D(D_4), .E(n6361), .C(wclk), .QN(n1604) );
  DFE1 \mem_reg_189][3  ( .D(D_3), .E(n6361), .C(wclk), .QN(n1605) );
  DFE1 \mem_reg_189][2  ( .D(D_2), .E(n6361), .C(wclk), .QN(n1606) );
  DFE1 \mem_reg_189][1  ( .D(D_1), .E(n6361), .C(wclk), .QN(n1607) );
  DFE1 \mem_reg_189][0  ( .D(D_0), .E(n6361), .C(wclk), .QN(n1608) );
  DFE1 \mem_reg_188][23  ( .D(D_23), .E(n6360), .C(wclk), .QN(n1609) );
  DFE1 \mem_reg_188][22  ( .D(D_22), .E(n6360), .C(wclk), .QN(n1610) );
  DFE1 \mem_reg_188][21  ( .D(D_21), .E(n6360), .C(wclk), .QN(n1611) );
  DFE1 \mem_reg_188][20  ( .D(D_20), .E(n6360), .C(wclk), .QN(n1612) );
  DFE1 \mem_reg_188][19  ( .D(D_19), .E(n6360), .C(wclk), .QN(n1613) );
  DFE1 \mem_reg_188][18  ( .D(D_18), .E(n6360), .C(wclk), .QN(n1614) );
  DFE1 \mem_reg_188][17  ( .D(D_17), .E(n6360), .C(wclk), .QN(n1615) );
  DFE1 \mem_reg_188][16  ( .D(D_16), .E(n6360), .C(wclk), .QN(n1616) );
  DFE1 \mem_reg_188][15  ( .D(D_15), .E(n6360), .C(wclk), .QN(n1617) );
  DFE1 \mem_reg_188][14  ( .D(D_14), .E(n6360), .C(wclk), .QN(n1618) );
  DFE1 \mem_reg_188][13  ( .D(D_13), .E(n6360), .C(wclk), .QN(n1619) );
  DFE1 \mem_reg_188][12  ( .D(D_12), .E(n6360), .C(wclk), .QN(n1620) );
  DFE1 \mem_reg_188][11  ( .D(D_11), .E(n6360), .C(wclk), .QN(n1621) );
  DFE1 \mem_reg_188][10  ( .D(D_10), .E(n6360), .C(wclk), .QN(n1622) );
  DFE1 \mem_reg_188][9  ( .D(D_9), .E(n6360), .C(wclk), .QN(n1623) );
  DFE1 \mem_reg_188][8  ( .D(D_8), .E(n6360), .C(wclk), .QN(n1624) );
  DFE1 \mem_reg_188][7  ( .D(D_7), .E(n6360), .C(wclk), .QN(n1625) );
  DFE1 \mem_reg_188][6  ( .D(D_6), .E(n6360), .C(wclk), .QN(n1626) );
  DFE1 \mem_reg_188][5  ( .D(D_5), .E(n6360), .C(wclk), .QN(n1627) );
  DFE1 \mem_reg_188][4  ( .D(D_4), .E(n6360), .C(wclk), .QN(n1628) );
  DFE1 \mem_reg_188][3  ( .D(D_3), .E(n6360), .C(wclk), .QN(n1629) );
  DFE1 \mem_reg_188][2  ( .D(D_2), .E(n6360), .C(wclk), .QN(n1630) );
  DFE1 \mem_reg_188][1  ( .D(D_1), .E(n6360), .C(wclk), .QN(n1631) );
  DFE1 \mem_reg_188][0  ( .D(D_0), .E(n6360), .C(wclk), .QN(n1632) );
  DFE1 \mem_reg_187][23  ( .D(D_23), .E(n6359), .C(wclk), .QN(n1633) );
  DFE1 \mem_reg_187][22  ( .D(D_22), .E(n6359), .C(wclk), .QN(n1634) );
  DFE1 \mem_reg_187][21  ( .D(D_21), .E(n6359), .C(wclk), .QN(n1635) );
  DFE1 \mem_reg_187][20  ( .D(D_20), .E(n6359), .C(wclk), .QN(n1636) );
  DFE1 \mem_reg_187][19  ( .D(D_19), .E(n6359), .C(wclk), .QN(n1637) );
  DFE1 \mem_reg_187][18  ( .D(D_18), .E(n6359), .C(wclk), .QN(n1638) );
  DFE1 \mem_reg_187][17  ( .D(D_17), .E(n6359), .C(wclk), .QN(n1639) );
  DFE1 \mem_reg_187][16  ( .D(D_16), .E(n6359), .C(wclk), .QN(n1640) );
  DFE1 \mem_reg_187][15  ( .D(D_15), .E(n6359), .C(wclk), .QN(n1641) );
  DFE1 \mem_reg_187][14  ( .D(D_14), .E(n6359), .C(wclk), .QN(n1642) );
  DFE1 \mem_reg_187][13  ( .D(D_13), .E(n6359), .C(wclk), .QN(n1643) );
  DFE1 \mem_reg_187][12  ( .D(D_12), .E(n6359), .C(wclk), .QN(n1644) );
  DFE1 \mem_reg_187][11  ( .D(D_11), .E(n6359), .C(wclk), .QN(n1645) );
  DFE1 \mem_reg_187][10  ( .D(D_10), .E(n6359), .C(wclk), .QN(n1646) );
  DFE1 \mem_reg_187][9  ( .D(D_9), .E(n6359), .C(wclk), .QN(n1647) );
  DFE1 \mem_reg_187][8  ( .D(D_8), .E(n6359), .C(wclk), .QN(n1648) );
  DFE1 \mem_reg_187][7  ( .D(D_7), .E(n6359), .C(wclk), .QN(n1649) );
  DFE1 \mem_reg_187][6  ( .D(D_6), .E(n6359), .C(wclk), .QN(n1650) );
  DFE1 \mem_reg_187][5  ( .D(D_5), .E(n6359), .C(wclk), .QN(n1651) );
  DFE1 \mem_reg_187][4  ( .D(D_4), .E(n6359), .C(wclk), .QN(n1652) );
  DFE1 \mem_reg_187][3  ( .D(D_3), .E(n6359), .C(wclk), .QN(n1653) );
  DFE1 \mem_reg_187][2  ( .D(D_2), .E(n6359), .C(wclk), .QN(n1654) );
  DFE1 \mem_reg_187][1  ( .D(D_1), .E(n6359), .C(wclk), .QN(n1655) );
  DFE1 \mem_reg_187][0  ( .D(D_0), .E(n6359), .C(wclk), .QN(n1656) );
  DFE1 \mem_reg_186][23  ( .D(D_23), .E(n6358), .C(wclk), .QN(n1657) );
  DFE1 \mem_reg_186][22  ( .D(D_22), .E(n6358), .C(wclk), .QN(n1658) );
  DFE1 \mem_reg_186][21  ( .D(D_21), .E(n6358), .C(wclk), .QN(n1659) );
  DFE1 \mem_reg_186][20  ( .D(D_20), .E(n6358), .C(wclk), .QN(n1660) );
  DFE1 \mem_reg_186][19  ( .D(D_19), .E(n6358), .C(wclk), .QN(n1661) );
  DFE1 \mem_reg_186][18  ( .D(D_18), .E(n6358), .C(wclk), .QN(n1662) );
  DFE1 \mem_reg_186][17  ( .D(D_17), .E(n6358), .C(wclk), .QN(n1663) );
  DFE1 \mem_reg_186][16  ( .D(D_16), .E(n6358), .C(wclk), .QN(n1664) );
  DFE1 \mem_reg_186][15  ( .D(D_15), .E(n6358), .C(wclk), .QN(n1665) );
  DFE1 \mem_reg_186][14  ( .D(D_14), .E(n6358), .C(wclk), .QN(n1666) );
  DFE1 \mem_reg_186][13  ( .D(D_13), .E(n6358), .C(wclk), .QN(n1667) );
  DFE1 \mem_reg_186][12  ( .D(D_12), .E(n6358), .C(wclk), .QN(n1668) );
  DFE1 \mem_reg_186][11  ( .D(D_11), .E(n6358), .C(wclk), .QN(n1669) );
  DFE1 \mem_reg_186][10  ( .D(D_10), .E(n6358), .C(wclk), .QN(n1670) );
  DFE1 \mem_reg_186][9  ( .D(D_9), .E(n6358), .C(wclk), .QN(n1671) );
  DFE1 \mem_reg_186][8  ( .D(D_8), .E(n6358), .C(wclk), .QN(n1672) );
  DFE1 \mem_reg_186][7  ( .D(D_7), .E(n6358), .C(wclk), .QN(n1673) );
  DFE1 \mem_reg_186][6  ( .D(D_6), .E(n6358), .C(wclk), .QN(n1674) );
  DFE1 \mem_reg_186][5  ( .D(D_5), .E(n6358), .C(wclk), .QN(n1675) );
  DFE1 \mem_reg_186][4  ( .D(D_4), .E(n6358), .C(wclk), .QN(n1676) );
  DFE1 \mem_reg_186][3  ( .D(D_3), .E(n6358), .C(wclk), .QN(n1677) );
  DFE1 \mem_reg_186][2  ( .D(D_2), .E(n6358), .C(wclk), .QN(n1678) );
  DFE1 \mem_reg_186][1  ( .D(D_1), .E(n6358), .C(wclk), .QN(n1679) );
  DFE1 \mem_reg_186][0  ( .D(D_0), .E(n6358), .C(wclk), .QN(n1680) );
  DFE1 \mem_reg_185][23  ( .D(D_23), .E(n6357), .C(wclk), .QN(n1681) );
  DFE1 \mem_reg_185][22  ( .D(D_22), .E(n6357), .C(wclk), .QN(n1682) );
  DFE1 \mem_reg_185][21  ( .D(D_21), .E(n6357), .C(wclk), .QN(n1683) );
  DFE1 \mem_reg_185][20  ( .D(D_20), .E(n6357), .C(wclk), .QN(n1684) );
  DFE1 \mem_reg_185][19  ( .D(D_19), .E(n6357), .C(wclk), .QN(n1685) );
  DFE1 \mem_reg_185][18  ( .D(D_18), .E(n6357), .C(wclk), .QN(n1686) );
  DFE1 \mem_reg_185][17  ( .D(D_17), .E(n6357), .C(wclk), .QN(n1687) );
  DFE1 \mem_reg_185][16  ( .D(D_16), .E(n6357), .C(wclk), .QN(n1688) );
  DFE1 \mem_reg_185][15  ( .D(D_15), .E(n6357), .C(wclk), .QN(n1689) );
  DFE1 \mem_reg_185][14  ( .D(D_14), .E(n6357), .C(wclk), .QN(n1690) );
  DFE1 \mem_reg_185][13  ( .D(D_13), .E(n6357), .C(wclk), .QN(n1691) );
  DFE1 \mem_reg_185][12  ( .D(D_12), .E(n6357), .C(wclk), .QN(n1692) );
  DFE1 \mem_reg_185][11  ( .D(D_11), .E(n6357), .C(wclk), .QN(n1693) );
  DFE1 \mem_reg_185][10  ( .D(D_10), .E(n6357), .C(wclk), .QN(n1694) );
  DFE1 \mem_reg_185][9  ( .D(D_9), .E(n6357), .C(wclk), .QN(n1695) );
  DFE1 \mem_reg_185][8  ( .D(D_8), .E(n6357), .C(wclk), .QN(n1696) );
  DFE1 \mem_reg_185][7  ( .D(D_7), .E(n6357), .C(wclk), .QN(n1697) );
  DFE1 \mem_reg_185][6  ( .D(D_6), .E(n6357), .C(wclk), .QN(n1698) );
  DFE1 \mem_reg_185][5  ( .D(D_5), .E(n6357), .C(wclk), .QN(n1699) );
  DFE1 \mem_reg_185][4  ( .D(D_4), .E(n6357), .C(wclk), .QN(n1700) );
  DFE1 \mem_reg_185][3  ( .D(D_3), .E(n6357), .C(wclk), .QN(n1701) );
  DFE1 \mem_reg_185][2  ( .D(D_2), .E(n6357), .C(wclk), .QN(n1702) );
  DFE1 \mem_reg_185][1  ( .D(D_1), .E(n6357), .C(wclk), .QN(n1703) );
  DFE1 \mem_reg_185][0  ( .D(D_0), .E(n6357), .C(wclk), .QN(n1704) );
  DFE1 \mem_reg_184][23  ( .D(D_23), .E(n6356), .C(wclk), .QN(n1705) );
  DFE1 \mem_reg_184][22  ( .D(D_22), .E(n6356), .C(wclk), .QN(n1706) );
  DFE1 \mem_reg_184][21  ( .D(D_21), .E(n6356), .C(wclk), .QN(n1707) );
  DFE1 \mem_reg_184][20  ( .D(D_20), .E(n6356), .C(wclk), .QN(n1708) );
  DFE1 \mem_reg_184][19  ( .D(D_19), .E(n6356), .C(wclk), .QN(n1709) );
  DFE1 \mem_reg_184][18  ( .D(D_18), .E(n6356), .C(wclk), .QN(n1710) );
  DFE1 \mem_reg_184][17  ( .D(D_17), .E(n6356), .C(wclk), .QN(n1711) );
  DFE1 \mem_reg_184][16  ( .D(D_16), .E(n6356), .C(wclk), .QN(n1712) );
  DFE1 \mem_reg_184][15  ( .D(D_15), .E(n6356), .C(wclk), .QN(n1713) );
  DFE1 \mem_reg_184][14  ( .D(D_14), .E(n6356), .C(wclk), .QN(n1714) );
  DFE1 \mem_reg_184][13  ( .D(D_13), .E(n6356), .C(wclk), .QN(n1715) );
  DFE1 \mem_reg_184][12  ( .D(D_12), .E(n6356), .C(wclk), .QN(n1716) );
  DFE1 \mem_reg_184][11  ( .D(D_11), .E(n6356), .C(wclk), .QN(n1717) );
  DFE1 \mem_reg_184][10  ( .D(D_10), .E(n6356), .C(wclk), .QN(n1718) );
  DFE1 \mem_reg_184][9  ( .D(D_9), .E(n6356), .C(wclk), .QN(n1719) );
  DFE1 \mem_reg_184][8  ( .D(D_8), .E(n6356), .C(wclk), .QN(n1720) );
  DFE1 \mem_reg_184][7  ( .D(D_7), .E(n6356), .C(wclk), .QN(n1721) );
  DFE1 \mem_reg_184][6  ( .D(D_6), .E(n6356), .C(wclk), .QN(n1722) );
  DFE1 \mem_reg_184][5  ( .D(D_5), .E(n6356), .C(wclk), .QN(n1723) );
  DFE1 \mem_reg_184][4  ( .D(D_4), .E(n6356), .C(wclk), .QN(n1724) );
  DFE1 \mem_reg_184][3  ( .D(D_3), .E(n6356), .C(wclk), .QN(n1725) );
  DFE1 \mem_reg_184][2  ( .D(D_2), .E(n6356), .C(wclk), .QN(n1726) );
  DFE1 \mem_reg_184][1  ( .D(D_1), .E(n6356), .C(wclk), .QN(n1727) );
  DFE1 \mem_reg_184][0  ( .D(D_0), .E(n6356), .C(wclk), .QN(n1728) );
  DFE1 \mem_reg_183][23  ( .D(D_23), .E(n6355), .C(wclk), .QN(n1729) );
  DFE1 \mem_reg_183][22  ( .D(D_22), .E(n6355), .C(wclk), .QN(n1730) );
  DFE1 \mem_reg_183][21  ( .D(D_21), .E(n6355), .C(wclk), .QN(n1731) );
  DFE1 \mem_reg_183][20  ( .D(D_20), .E(n6355), .C(wclk), .QN(n1732) );
  DFE1 \mem_reg_183][19  ( .D(D_19), .E(n6355), .C(wclk), .QN(n1733) );
  DFE1 \mem_reg_183][18  ( .D(D_18), .E(n6355), .C(wclk), .QN(n1734) );
  DFE1 \mem_reg_183][17  ( .D(D_17), .E(n6355), .C(wclk), .QN(n1735) );
  DFE1 \mem_reg_183][16  ( .D(D_16), .E(n6355), .C(wclk), .QN(n1736) );
  DFE1 \mem_reg_183][15  ( .D(D_15), .E(n6355), .C(wclk), .QN(n1737) );
  DFE1 \mem_reg_183][14  ( .D(D_14), .E(n6355), .C(wclk), .QN(n1738) );
  DFE1 \mem_reg_183][13  ( .D(D_13), .E(n6355), .C(wclk), .QN(n1739) );
  DFE1 \mem_reg_183][12  ( .D(D_12), .E(n6355), .C(wclk), .QN(n1740) );
  DFE1 \mem_reg_183][11  ( .D(D_11), .E(n6355), .C(wclk), .QN(n1741) );
  DFE1 \mem_reg_183][10  ( .D(D_10), .E(n6355), .C(wclk), .QN(n1742) );
  DFE1 \mem_reg_183][9  ( .D(D_9), .E(n6355), .C(wclk), .QN(n1743) );
  DFE1 \mem_reg_183][8  ( .D(D_8), .E(n6355), .C(wclk), .QN(n1744) );
  DFE1 \mem_reg_183][7  ( .D(D_7), .E(n6355), .C(wclk), .QN(n1745) );
  DFE1 \mem_reg_183][6  ( .D(D_6), .E(n6355), .C(wclk), .QN(n1746) );
  DFE1 \mem_reg_183][5  ( .D(D_5), .E(n6355), .C(wclk), .QN(n1747) );
  DFE1 \mem_reg_183][4  ( .D(D_4), .E(n6355), .C(wclk), .QN(n1748) );
  DFE1 \mem_reg_183][3  ( .D(D_3), .E(n6355), .C(wclk), .QN(n1749) );
  DFE1 \mem_reg_183][2  ( .D(D_2), .E(n6355), .C(wclk), .QN(n1750) );
  DFE1 \mem_reg_183][1  ( .D(D_1), .E(n6355), .C(wclk), .QN(n1751) );
  DFE1 \mem_reg_183][0  ( .D(D_0), .E(n6355), .C(wclk), .QN(n1752) );
  DFE1 \mem_reg_182][23  ( .D(D_23), .E(n6354), .C(wclk), .QN(n1753) );
  DFE1 \mem_reg_182][22  ( .D(D_22), .E(n6354), .C(wclk), .QN(n1754) );
  DFE1 \mem_reg_182][21  ( .D(D_21), .E(n6354), .C(wclk), .QN(n1755) );
  DFE1 \mem_reg_182][20  ( .D(D_20), .E(n6354), .C(wclk), .QN(n1756) );
  DFE1 \mem_reg_182][19  ( .D(D_19), .E(n6354), .C(wclk), .QN(n1757) );
  DFE1 \mem_reg_182][18  ( .D(D_18), .E(n6354), .C(wclk), .QN(n1758) );
  DFE1 \mem_reg_182][17  ( .D(D_17), .E(n6354), .C(wclk), .QN(n1759) );
  DFE1 \mem_reg_182][16  ( .D(D_16), .E(n6354), .C(wclk), .QN(n1760) );
  DFE1 \mem_reg_182][15  ( .D(D_15), .E(n6354), .C(wclk), .QN(n1761) );
  DFE1 \mem_reg_182][14  ( .D(D_14), .E(n6354), .C(wclk), .QN(n1762) );
  DFE1 \mem_reg_182][13  ( .D(D_13), .E(n6354), .C(wclk), .QN(n1763) );
  DFE1 \mem_reg_182][12  ( .D(D_12), .E(n6354), .C(wclk), .QN(n1764) );
  DFE1 \mem_reg_182][11  ( .D(D_11), .E(n6354), .C(wclk), .QN(n1765) );
  DFE1 \mem_reg_182][10  ( .D(D_10), .E(n6354), .C(wclk), .QN(n1766) );
  DFE1 \mem_reg_182][9  ( .D(D_9), .E(n6354), .C(wclk), .QN(n1767) );
  DFE1 \mem_reg_182][8  ( .D(D_8), .E(n6354), .C(wclk), .QN(n1768) );
  DFE1 \mem_reg_182][7  ( .D(D_7), .E(n6354), .C(wclk), .QN(n1769) );
  DFE1 \mem_reg_182][6  ( .D(D_6), .E(n6354), .C(wclk), .QN(n1770) );
  DFE1 \mem_reg_182][5  ( .D(D_5), .E(n6354), .C(wclk), .QN(n1771) );
  DFE1 \mem_reg_182][4  ( .D(D_4), .E(n6354), .C(wclk), .QN(n1772) );
  DFE1 \mem_reg_182][3  ( .D(D_3), .E(n6354), .C(wclk), .QN(n1773) );
  DFE1 \mem_reg_182][2  ( .D(D_2), .E(n6354), .C(wclk), .QN(n1774) );
  DFE1 \mem_reg_182][1  ( .D(D_1), .E(n6354), .C(wclk), .QN(n1775) );
  DFE1 \mem_reg_182][0  ( .D(D_0), .E(n6354), .C(wclk), .QN(n1776) );
  DFE1 \mem_reg_181][23  ( .D(D_23), .E(n6353), .C(wclk), .QN(n1777) );
  DFE1 \mem_reg_181][22  ( .D(D_22), .E(n6353), .C(wclk), .QN(n1778) );
  DFE1 \mem_reg_181][21  ( .D(D_21), .E(n6353), .C(wclk), .QN(n1779) );
  DFE1 \mem_reg_181][20  ( .D(D_20), .E(n6353), .C(wclk), .QN(n1780) );
  DFE1 \mem_reg_181][19  ( .D(D_19), .E(n6353), .C(wclk), .QN(n1781) );
  DFE1 \mem_reg_181][18  ( .D(D_18), .E(n6353), .C(wclk), .QN(n1782) );
  DFE1 \mem_reg_181][17  ( .D(D_17), .E(n6353), .C(wclk), .QN(n1783) );
  DFE1 \mem_reg_181][16  ( .D(D_16), .E(n6353), .C(wclk), .QN(n1784) );
  DFE1 \mem_reg_181][15  ( .D(D_15), .E(n6353), .C(wclk), .QN(n1785) );
  DFE1 \mem_reg_181][14  ( .D(D_14), .E(n6353), .C(wclk), .QN(n1786) );
  DFE1 \mem_reg_181][13  ( .D(D_13), .E(n6353), .C(wclk), .QN(n1787) );
  DFE1 \mem_reg_181][12  ( .D(D_12), .E(n6353), .C(wclk), .QN(n1788) );
  DFE1 \mem_reg_181][11  ( .D(D_11), .E(n6353), .C(wclk), .QN(n1789) );
  DFE1 \mem_reg_181][10  ( .D(D_10), .E(n6353), .C(wclk), .QN(n1790) );
  DFE1 \mem_reg_181][9  ( .D(D_9), .E(n6353), .C(wclk), .QN(n1791) );
  DFE1 \mem_reg_181][8  ( .D(D_8), .E(n6353), .C(wclk), .QN(n1792) );
  DFE1 \mem_reg_181][7  ( .D(D_7), .E(n6353), .C(wclk), .QN(n1793) );
  DFE1 \mem_reg_181][6  ( .D(D_6), .E(n6353), .C(wclk), .QN(n1794) );
  DFE1 \mem_reg_181][5  ( .D(D_5), .E(n6353), .C(wclk), .QN(n1795) );
  DFE1 \mem_reg_181][4  ( .D(D_4), .E(n6353), .C(wclk), .QN(n1796) );
  DFE1 \mem_reg_181][3  ( .D(D_3), .E(n6353), .C(wclk), .QN(n1797) );
  DFE1 \mem_reg_181][2  ( .D(D_2), .E(n6353), .C(wclk), .QN(n1798) );
  DFE1 \mem_reg_181][1  ( .D(D_1), .E(n6353), .C(wclk), .QN(n1799) );
  DFE1 \mem_reg_181][0  ( .D(D_0), .E(n6353), .C(wclk), .QN(n1800) );
  DFE1 \mem_reg_180][23  ( .D(D_23), .E(n6352), .C(wclk), .QN(n1801) );
  DFE1 \mem_reg_180][22  ( .D(D_22), .E(n6352), .C(wclk), .QN(n1802) );
  DFE1 \mem_reg_180][21  ( .D(D_21), .E(n6352), .C(wclk), .QN(n1803) );
  DFE1 \mem_reg_180][20  ( .D(D_20), .E(n6352), .C(wclk), .QN(n1804) );
  DFE1 \mem_reg_180][19  ( .D(D_19), .E(n6352), .C(wclk), .QN(n1805) );
  DFE1 \mem_reg_180][18  ( .D(D_18), .E(n6352), .C(wclk), .QN(n1806) );
  DFE1 \mem_reg_180][17  ( .D(D_17), .E(n6352), .C(wclk), .QN(n1807) );
  DFE1 \mem_reg_180][16  ( .D(D_16), .E(n6352), .C(wclk), .QN(n1808) );
  DFE1 \mem_reg_180][15  ( .D(D_15), .E(n6352), .C(wclk), .QN(n1809) );
  DFE1 \mem_reg_180][14  ( .D(D_14), .E(n6352), .C(wclk), .QN(n1810) );
  DFE1 \mem_reg_180][13  ( .D(D_13), .E(n6352), .C(wclk), .QN(n1811) );
  DFE1 \mem_reg_180][12  ( .D(D_12), .E(n6352), .C(wclk), .QN(n1812) );
  DFE1 \mem_reg_180][11  ( .D(D_11), .E(n6352), .C(wclk), .QN(n1813) );
  DFE1 \mem_reg_180][10  ( .D(D_10), .E(n6352), .C(wclk), .QN(n1814) );
  DFE1 \mem_reg_180][9  ( .D(D_9), .E(n6352), .C(wclk), .QN(n1815) );
  DFE1 \mem_reg_180][8  ( .D(D_8), .E(n6352), .C(wclk), .QN(n1816) );
  DFE1 \mem_reg_180][7  ( .D(D_7), .E(n6352), .C(wclk), .QN(n1817) );
  DFE1 \mem_reg_180][6  ( .D(D_6), .E(n6352), .C(wclk), .QN(n1818) );
  DFE1 \mem_reg_180][5  ( .D(D_5), .E(n6352), .C(wclk), .QN(n1819) );
  DFE1 \mem_reg_180][4  ( .D(D_4), .E(n6352), .C(wclk), .QN(n1820) );
  DFE1 \mem_reg_180][3  ( .D(D_3), .E(n6352), .C(wclk), .QN(n1821) );
  DFE1 \mem_reg_180][2  ( .D(D_2), .E(n6352), .C(wclk), .QN(n1822) );
  DFE1 \mem_reg_180][1  ( .D(D_1), .E(n6352), .C(wclk), .QN(n1823) );
  DFE1 \mem_reg_180][0  ( .D(D_0), .E(n6352), .C(wclk), .QN(n1824) );
  DFE1 \mem_reg_179][23  ( .D(D_23), .E(n6351), .C(wclk), .QN(n1825) );
  DFE1 \mem_reg_179][22  ( .D(D_22), .E(n6351), .C(wclk), .QN(n1826) );
  DFE1 \mem_reg_179][21  ( .D(D_21), .E(n6351), .C(wclk), .QN(n1827) );
  DFE1 \mem_reg_179][20  ( .D(D_20), .E(n6351), .C(wclk), .QN(n1828) );
  DFE1 \mem_reg_179][19  ( .D(D_19), .E(n6351), .C(wclk), .QN(n1829) );
  DFE1 \mem_reg_179][18  ( .D(D_18), .E(n6351), .C(wclk), .QN(n1830) );
  DFE1 \mem_reg_179][17  ( .D(D_17), .E(n6351), .C(wclk), .QN(n1831) );
  DFE1 \mem_reg_179][16  ( .D(D_16), .E(n6351), .C(wclk), .QN(n1832) );
  DFE1 \mem_reg_179][15  ( .D(D_15), .E(n6351), .C(wclk), .QN(n1833) );
  DFE1 \mem_reg_179][14  ( .D(D_14), .E(n6351), .C(wclk), .QN(n1834) );
  DFE1 \mem_reg_179][13  ( .D(D_13), .E(n6351), .C(wclk), .QN(n1835) );
  DFE1 \mem_reg_179][12  ( .D(D_12), .E(n6351), .C(wclk), .QN(n1836) );
  DFE1 \mem_reg_179][11  ( .D(D_11), .E(n6351), .C(wclk), .QN(n1837) );
  DFE1 \mem_reg_179][10  ( .D(D_10), .E(n6351), .C(wclk), .QN(n1838) );
  DFE1 \mem_reg_179][9  ( .D(D_9), .E(n6351), .C(wclk), .QN(n1839) );
  DFE1 \mem_reg_179][8  ( .D(D_8), .E(n6351), .C(wclk), .QN(n1840) );
  DFE1 \mem_reg_179][7  ( .D(D_7), .E(n6351), .C(wclk), .QN(n1841) );
  DFE1 \mem_reg_179][6  ( .D(D_6), .E(n6351), .C(wclk), .QN(n1842) );
  DFE1 \mem_reg_179][5  ( .D(D_5), .E(n6351), .C(wclk), .QN(n1843) );
  DFE1 \mem_reg_179][4  ( .D(D_4), .E(n6351), .C(wclk), .QN(n1844) );
  DFE1 \mem_reg_179][3  ( .D(D_3), .E(n6351), .C(wclk), .QN(n1845) );
  DFE1 \mem_reg_179][2  ( .D(D_2), .E(n6351), .C(wclk), .QN(n1846) );
  DFE1 \mem_reg_179][1  ( .D(D_1), .E(n6351), .C(wclk), .QN(n1847) );
  DFE1 \mem_reg_179][0  ( .D(D_0), .E(n6351), .C(wclk), .QN(n1848) );
  DFE1 \mem_reg_178][23  ( .D(D_23), .E(n6350), .C(wclk), .QN(n1849) );
  DFE1 \mem_reg_178][22  ( .D(D_22), .E(n6350), .C(wclk), .QN(n1850) );
  DFE1 \mem_reg_178][21  ( .D(D_21), .E(n6350), .C(wclk), .QN(n1851) );
  DFE1 \mem_reg_178][20  ( .D(D_20), .E(n6350), .C(wclk), .QN(n1852) );
  DFE1 \mem_reg_178][19  ( .D(D_19), .E(n6350), .C(wclk), .QN(n1853) );
  DFE1 \mem_reg_178][18  ( .D(D_18), .E(n6350), .C(wclk), .QN(n1854) );
  DFE1 \mem_reg_178][17  ( .D(D_17), .E(n6350), .C(wclk), .QN(n1855) );
  DFE1 \mem_reg_178][16  ( .D(D_16), .E(n6350), .C(wclk), .QN(n1856) );
  DFE1 \mem_reg_178][15  ( .D(D_15), .E(n6350), .C(wclk), .QN(n1857) );
  DFE1 \mem_reg_178][14  ( .D(D_14), .E(n6350), .C(wclk), .QN(n1858) );
  DFE1 \mem_reg_178][13  ( .D(D_13), .E(n6350), .C(wclk), .QN(n1859) );
  DFE1 \mem_reg_178][12  ( .D(D_12), .E(n6350), .C(wclk), .QN(n1860) );
  DFE1 \mem_reg_178][11  ( .D(D_11), .E(n6350), .C(wclk), .QN(n1861) );
  DFE1 \mem_reg_178][10  ( .D(D_10), .E(n6350), .C(wclk), .QN(n1862) );
  DFE1 \mem_reg_178][9  ( .D(D_9), .E(n6350), .C(wclk), .QN(n1863) );
  DFE1 \mem_reg_178][8  ( .D(D_8), .E(n6350), .C(wclk), .QN(n1864) );
  DFE1 \mem_reg_178][7  ( .D(D_7), .E(n6350), .C(wclk), .QN(n1865) );
  DFE1 \mem_reg_178][6  ( .D(D_6), .E(n6350), .C(wclk), .QN(n1866) );
  DFE1 \mem_reg_178][5  ( .D(D_5), .E(n6350), .C(wclk), .QN(n1867) );
  DFE1 \mem_reg_178][4  ( .D(D_4), .E(n6350), .C(wclk), .QN(n1868) );
  DFE1 \mem_reg_178][3  ( .D(D_3), .E(n6350), .C(wclk), .QN(n1869) );
  DFE1 \mem_reg_178][2  ( .D(D_2), .E(n6350), .C(wclk), .QN(n1870) );
  DFE1 \mem_reg_178][1  ( .D(D_1), .E(n6350), .C(wclk), .QN(n1871) );
  DFE1 \mem_reg_178][0  ( .D(D_0), .E(n6350), .C(wclk), .QN(n1872) );
  DFE1 \mem_reg_177][23  ( .D(D_23), .E(n6349), .C(wclk), .QN(n1873) );
  DFE1 \mem_reg_177][22  ( .D(D_22), .E(n6349), .C(wclk), .QN(n1874) );
  DFE1 \mem_reg_177][21  ( .D(D_21), .E(n6349), .C(wclk), .QN(n1875) );
  DFE1 \mem_reg_177][20  ( .D(D_20), .E(n6349), .C(wclk), .QN(n1876) );
  DFE1 \mem_reg_177][19  ( .D(D_19), .E(n6349), .C(wclk), .QN(n1877) );
  DFE1 \mem_reg_177][18  ( .D(D_18), .E(n6349), .C(wclk), .QN(n1878) );
  DFE1 \mem_reg_177][17  ( .D(D_17), .E(n6349), .C(wclk), .QN(n1879) );
  DFE1 \mem_reg_177][16  ( .D(D_16), .E(n6349), .C(wclk), .QN(n1880) );
  DFE1 \mem_reg_177][15  ( .D(D_15), .E(n6349), .C(wclk), .QN(n1881) );
  DFE1 \mem_reg_177][14  ( .D(D_14), .E(n6349), .C(wclk), .QN(n1882) );
  DFE1 \mem_reg_177][13  ( .D(D_13), .E(n6349), .C(wclk), .QN(n1883) );
  DFE1 \mem_reg_177][12  ( .D(D_12), .E(n6349), .C(wclk), .QN(n1884) );
  DFE1 \mem_reg_177][11  ( .D(D_11), .E(n6349), .C(wclk), .QN(n1885) );
  DFE1 \mem_reg_177][10  ( .D(D_10), .E(n6349), .C(wclk), .QN(n1886) );
  DFE1 \mem_reg_177][9  ( .D(D_9), .E(n6349), .C(wclk), .QN(n1887) );
  DFE1 \mem_reg_177][8  ( .D(D_8), .E(n6349), .C(wclk), .QN(n1888) );
  DFE1 \mem_reg_177][7  ( .D(D_7), .E(n6349), .C(wclk), .QN(n1889) );
  DFE1 \mem_reg_177][6  ( .D(D_6), .E(n6349), .C(wclk), .QN(n1890) );
  DFE1 \mem_reg_177][5  ( .D(D_5), .E(n6349), .C(wclk), .QN(n1891) );
  DFE1 \mem_reg_177][4  ( .D(D_4), .E(n6349), .C(wclk), .QN(n1892) );
  DFE1 \mem_reg_177][3  ( .D(D_3), .E(n6349), .C(wclk), .QN(n1893) );
  DFE1 \mem_reg_177][2  ( .D(D_2), .E(n6349), .C(wclk), .QN(n1894) );
  DFE1 \mem_reg_177][1  ( .D(D_1), .E(n6349), .C(wclk), .QN(n1895) );
  DFE1 \mem_reg_177][0  ( .D(D_0), .E(n6349), .C(wclk), .QN(n1896) );
  DFE1 \mem_reg_176][23  ( .D(D_23), .E(n6347), .C(wclk), .QN(n1897) );
  DFE1 \mem_reg_176][22  ( .D(D_22), .E(n6347), .C(wclk), .QN(n1898) );
  DFE1 \mem_reg_176][21  ( .D(D_21), .E(n6347), .C(wclk), .QN(n1899) );
  DFE1 \mem_reg_176][20  ( .D(D_20), .E(n6347), .C(wclk), .QN(n1900) );
  DFE1 \mem_reg_176][19  ( .D(D_19), .E(n6347), .C(wclk), .QN(n1901) );
  DFE1 \mem_reg_176][18  ( .D(D_18), .E(n6347), .C(wclk), .QN(n1902) );
  DFE1 \mem_reg_176][17  ( .D(D_17), .E(n6347), .C(wclk), .QN(n1903) );
  DFE1 \mem_reg_176][16  ( .D(D_16), .E(n6347), .C(wclk), .QN(n1904) );
  DFE1 \mem_reg_176][15  ( .D(D_15), .E(n6347), .C(wclk), .QN(n1905) );
  DFE1 \mem_reg_176][14  ( .D(D_14), .E(n6347), .C(wclk), .QN(n1906) );
  DFE1 \mem_reg_176][13  ( .D(D_13), .E(n6347), .C(wclk), .QN(n1907) );
  DFE1 \mem_reg_176][12  ( .D(D_12), .E(n6347), .C(wclk), .QN(n1908) );
  DFE1 \mem_reg_176][11  ( .D(D_11), .E(n6347), .C(wclk), .QN(n1909) );
  DFE1 \mem_reg_176][10  ( .D(D_10), .E(n6347), .C(wclk), .QN(n1910) );
  DFE1 \mem_reg_176][9  ( .D(D_9), .E(n6347), .C(wclk), .QN(n1911) );
  DFE1 \mem_reg_176][8  ( .D(D_8), .E(n6347), .C(wclk), .QN(n1912) );
  DFE1 \mem_reg_176][7  ( .D(D_7), .E(n6347), .C(wclk), .QN(n1913) );
  DFE1 \mem_reg_176][6  ( .D(D_6), .E(n6347), .C(wclk), .QN(n1914) );
  DFE1 \mem_reg_176][5  ( .D(D_5), .E(n6347), .C(wclk), .QN(n1915) );
  DFE1 \mem_reg_176][4  ( .D(D_4), .E(n6347), .C(wclk), .QN(n1916) );
  DFE1 \mem_reg_176][3  ( .D(D_3), .E(n6347), .C(wclk), .QN(n1917) );
  DFE1 \mem_reg_176][2  ( .D(D_2), .E(n6347), .C(wclk), .QN(n1918) );
  DFE1 \mem_reg_176][1  ( .D(D_1), .E(n6347), .C(wclk), .QN(n1919) );
  DFE1 \mem_reg_176][0  ( .D(D_0), .E(n6347), .C(wclk), .QN(n1920) );
  DFE1 \mem_reg_175][23  ( .D(D_23), .E(n6346), .C(wclk), .QN(n1921) );
  DFE1 \mem_reg_175][22  ( .D(D_22), .E(n6346), .C(wclk), .QN(n1922) );
  DFE1 \mem_reg_175][21  ( .D(D_21), .E(n6346), .C(wclk), .QN(n1923) );
  DFE1 \mem_reg_175][20  ( .D(D_20), .E(n6346), .C(wclk), .QN(n1924) );
  DFE1 \mem_reg_175][19  ( .D(D_19), .E(n6346), .C(wclk), .QN(n1925) );
  DFE1 \mem_reg_175][18  ( .D(D_18), .E(n6346), .C(wclk), .QN(n1926) );
  DFE1 \mem_reg_175][17  ( .D(D_17), .E(n6346), .C(wclk), .QN(n1927) );
  DFE1 \mem_reg_175][16  ( .D(D_16), .E(n6346), .C(wclk), .QN(n1928) );
  DFE1 \mem_reg_175][15  ( .D(D_15), .E(n6346), .C(wclk), .QN(n1929) );
  DFE1 \mem_reg_175][14  ( .D(D_14), .E(n6346), .C(wclk), .QN(n1930) );
  DFE1 \mem_reg_175][13  ( .D(D_13), .E(n6346), .C(wclk), .QN(n1931) );
  DFE1 \mem_reg_175][12  ( .D(D_12), .E(n6346), .C(wclk), .QN(n1932) );
  DFE1 \mem_reg_175][11  ( .D(D_11), .E(n6346), .C(wclk), .QN(n1933) );
  DFE1 \mem_reg_175][10  ( .D(D_10), .E(n6346), .C(wclk), .QN(n1934) );
  DFE1 \mem_reg_175][9  ( .D(D_9), .E(n6346), .C(wclk), .QN(n1935) );
  DFE1 \mem_reg_175][8  ( .D(D_8), .E(n6346), .C(wclk), .QN(n1936) );
  DFE1 \mem_reg_175][7  ( .D(D_7), .E(n6346), .C(wclk), .QN(n1937) );
  DFE1 \mem_reg_175][6  ( .D(D_6), .E(n6346), .C(wclk), .QN(n1938) );
  DFE1 \mem_reg_175][5  ( .D(D_5), .E(n6346), .C(wclk), .QN(n1939) );
  DFE1 \mem_reg_175][4  ( .D(D_4), .E(n6346), .C(wclk), .QN(n1940) );
  DFE1 \mem_reg_175][3  ( .D(D_3), .E(n6346), .C(wclk), .QN(n1941) );
  DFE1 \mem_reg_175][2  ( .D(D_2), .E(n6346), .C(wclk), .QN(n1942) );
  DFE1 \mem_reg_175][1  ( .D(D_1), .E(n6346), .C(wclk), .QN(n1943) );
  DFE1 \mem_reg_175][0  ( .D(D_0), .E(n6346), .C(wclk), .QN(n1944) );
  DFE1 \mem_reg_174][23  ( .D(D_23), .E(n6345), .C(wclk), .QN(n1945) );
  DFE1 \mem_reg_174][22  ( .D(D_22), .E(n6345), .C(wclk), .QN(n1946) );
  DFE1 \mem_reg_174][21  ( .D(D_21), .E(n6345), .C(wclk), .QN(n1947) );
  DFE1 \mem_reg_174][20  ( .D(D_20), .E(n6345), .C(wclk), .QN(n1948) );
  DFE1 \mem_reg_174][19  ( .D(D_19), .E(n6345), .C(wclk), .QN(n1949) );
  DFE1 \mem_reg_174][18  ( .D(D_18), .E(n6345), .C(wclk), .QN(n1950) );
  DFE1 \mem_reg_174][17  ( .D(D_17), .E(n6345), .C(wclk), .QN(n1951) );
  DFE1 \mem_reg_174][16  ( .D(D_16), .E(n6345), .C(wclk), .QN(n1952) );
  DFE1 \mem_reg_174][15  ( .D(D_15), .E(n6345), .C(wclk), .QN(n1953) );
  DFE1 \mem_reg_174][14  ( .D(D_14), .E(n6345), .C(wclk), .QN(n1954) );
  DFE1 \mem_reg_174][13  ( .D(D_13), .E(n6345), .C(wclk), .QN(n1955) );
  DFE1 \mem_reg_174][12  ( .D(D_12), .E(n6345), .C(wclk), .QN(n1956) );
  DFE1 \mem_reg_174][11  ( .D(D_11), .E(n6345), .C(wclk), .QN(n1957) );
  DFE1 \mem_reg_174][10  ( .D(D_10), .E(n6345), .C(wclk), .QN(n1958) );
  DFE1 \mem_reg_174][9  ( .D(D_9), .E(n6345), .C(wclk), .QN(n1959) );
  DFE1 \mem_reg_174][8  ( .D(D_8), .E(n6345), .C(wclk), .QN(n1960) );
  DFE1 \mem_reg_174][7  ( .D(D_7), .E(n6345), .C(wclk), .QN(n1961) );
  DFE1 \mem_reg_174][6  ( .D(D_6), .E(n6345), .C(wclk), .QN(n1962) );
  DFE1 \mem_reg_174][5  ( .D(D_5), .E(n6345), .C(wclk), .QN(n1963) );
  DFE1 \mem_reg_174][4  ( .D(D_4), .E(n6345), .C(wclk), .QN(n1964) );
  DFE1 \mem_reg_174][3  ( .D(D_3), .E(n6345), .C(wclk), .QN(n1965) );
  DFE1 \mem_reg_174][2  ( .D(D_2), .E(n6345), .C(wclk), .QN(n1966) );
  DFE1 \mem_reg_174][1  ( .D(D_1), .E(n6345), .C(wclk), .QN(n1967) );
  DFE1 \mem_reg_174][0  ( .D(D_0), .E(n6345), .C(wclk), .QN(n1968) );
  DFE1 \mem_reg_173][23  ( .D(D_23), .E(n6344), .C(wclk), .QN(n1969) );
  DFE1 \mem_reg_173][22  ( .D(D_22), .E(n6344), .C(wclk), .QN(n1970) );
  DFE1 \mem_reg_173][21  ( .D(D_21), .E(n6344), .C(wclk), .QN(n1971) );
  DFE1 \mem_reg_173][20  ( .D(D_20), .E(n6344), .C(wclk), .QN(n1972) );
  DFE1 \mem_reg_173][19  ( .D(D_19), .E(n6344), .C(wclk), .QN(n1973) );
  DFE1 \mem_reg_173][18  ( .D(D_18), .E(n6344), .C(wclk), .QN(n1974) );
  DFE1 \mem_reg_173][17  ( .D(D_17), .E(n6344), .C(wclk), .QN(n1975) );
  DFE1 \mem_reg_173][16  ( .D(D_16), .E(n6344), .C(wclk), .QN(n1976) );
  DFE1 \mem_reg_173][15  ( .D(D_15), .E(n6344), .C(wclk), .QN(n1977) );
  DFE1 \mem_reg_173][14  ( .D(D_14), .E(n6344), .C(wclk), .QN(n1978) );
  DFE1 \mem_reg_173][13  ( .D(D_13), .E(n6344), .C(wclk), .QN(n1979) );
  DFE1 \mem_reg_173][12  ( .D(D_12), .E(n6344), .C(wclk), .QN(n1980) );
  DFE1 \mem_reg_173][11  ( .D(D_11), .E(n6344), .C(wclk), .QN(n1981) );
  DFE1 \mem_reg_173][10  ( .D(D_10), .E(n6344), .C(wclk), .QN(n1982) );
  DFE1 \mem_reg_173][9  ( .D(D_9), .E(n6344), .C(wclk), .QN(n1983) );
  DFE1 \mem_reg_173][8  ( .D(D_8), .E(n6344), .C(wclk), .QN(n1984) );
  DFE1 \mem_reg_173][7  ( .D(D_7), .E(n6344), .C(wclk), .QN(n1985) );
  DFE1 \mem_reg_173][6  ( .D(D_6), .E(n6344), .C(wclk), .QN(n1986) );
  DFE1 \mem_reg_173][5  ( .D(D_5), .E(n6344), .C(wclk), .QN(n1987) );
  DFE1 \mem_reg_173][4  ( .D(D_4), .E(n6344), .C(wclk), .QN(n1988) );
  DFE1 \mem_reg_173][3  ( .D(D_3), .E(n6344), .C(wclk), .QN(n1989) );
  DFE1 \mem_reg_173][2  ( .D(D_2), .E(n6344), .C(wclk), .QN(n1990) );
  DFE1 \mem_reg_173][1  ( .D(D_1), .E(n6344), .C(wclk), .QN(n1991) );
  DFE1 \mem_reg_173][0  ( .D(D_0), .E(n6344), .C(wclk), .QN(n1992) );
  DFE1 \mem_reg_172][23  ( .D(D_23), .E(n6343), .C(wclk), .QN(n1993) );
  DFE1 \mem_reg_172][22  ( .D(D_22), .E(n6343), .C(wclk), .QN(n1994) );
  DFE1 \mem_reg_172][21  ( .D(D_21), .E(n6343), .C(wclk), .QN(n1995) );
  DFE1 \mem_reg_172][20  ( .D(D_20), .E(n6343), .C(wclk), .QN(n1996) );
  DFE1 \mem_reg_172][19  ( .D(D_19), .E(n6343), .C(wclk), .QN(n1997) );
  DFE1 \mem_reg_172][18  ( .D(D_18), .E(n6343), .C(wclk), .QN(n1998) );
  DFE1 \mem_reg_172][17  ( .D(D_17), .E(n6343), .C(wclk), .QN(n1999) );
  DFE1 \mem_reg_172][16  ( .D(D_16), .E(n6343), .C(wclk), .QN(n2000) );
  DFE1 \mem_reg_172][15  ( .D(D_15), .E(n6343), .C(wclk), .QN(n2001) );
  DFE1 \mem_reg_172][14  ( .D(D_14), .E(n6343), .C(wclk), .QN(n2002) );
  DFE1 \mem_reg_172][13  ( .D(D_13), .E(n6343), .C(wclk), .QN(n2003) );
  DFE1 \mem_reg_172][12  ( .D(D_12), .E(n6343), .C(wclk), .QN(n2004) );
  DFE1 \mem_reg_172][11  ( .D(D_11), .E(n6343), .C(wclk), .QN(n2005) );
  DFE1 \mem_reg_172][10  ( .D(D_10), .E(n6343), .C(wclk), .QN(n2006) );
  DFE1 \mem_reg_172][9  ( .D(D_9), .E(n6343), .C(wclk), .QN(n2007) );
  DFE1 \mem_reg_172][8  ( .D(D_8), .E(n6343), .C(wclk), .QN(n2008) );
  DFE1 \mem_reg_172][7  ( .D(D_7), .E(n6343), .C(wclk), .QN(n2009) );
  DFE1 \mem_reg_172][6  ( .D(D_6), .E(n6343), .C(wclk), .QN(n2010) );
  DFE1 \mem_reg_172][5  ( .D(D_5), .E(n6343), .C(wclk), .QN(n2011) );
  DFE1 \mem_reg_172][4  ( .D(D_4), .E(n6343), .C(wclk), .QN(n2012) );
  DFE1 \mem_reg_172][3  ( .D(D_3), .E(n6343), .C(wclk), .QN(n2013) );
  DFE1 \mem_reg_172][2  ( .D(D_2), .E(n6343), .C(wclk), .QN(n2014) );
  DFE1 \mem_reg_172][1  ( .D(D_1), .E(n6343), .C(wclk), .QN(n2015) );
  DFE1 \mem_reg_172][0  ( .D(D_0), .E(n6343), .C(wclk), .QN(n2016) );
  DFE1 \mem_reg_171][23  ( .D(D_23), .E(n6342), .C(wclk), .QN(n2017) );
  DFE1 \mem_reg_171][22  ( .D(D_22), .E(n6342), .C(wclk), .QN(n2018) );
  DFE1 \mem_reg_171][21  ( .D(D_21), .E(n6342), .C(wclk), .QN(n2019) );
  DFE1 \mem_reg_171][20  ( .D(D_20), .E(n6342), .C(wclk), .QN(n2020) );
  DFE1 \mem_reg_171][19  ( .D(D_19), .E(n6342), .C(wclk), .QN(n2021) );
  DFE1 \mem_reg_171][18  ( .D(D_18), .E(n6342), .C(wclk), .QN(n2022) );
  DFE1 \mem_reg_171][17  ( .D(D_17), .E(n6342), .C(wclk), .QN(n2023) );
  DFE1 \mem_reg_171][16  ( .D(D_16), .E(n6342), .C(wclk), .QN(n2024) );
  DFE1 \mem_reg_171][15  ( .D(D_15), .E(n6342), .C(wclk), .QN(n2025) );
  DFE1 \mem_reg_171][14  ( .D(D_14), .E(n6342), .C(wclk), .QN(n2026) );
  DFE1 \mem_reg_171][13  ( .D(D_13), .E(n6342), .C(wclk), .QN(n2027) );
  DFE1 \mem_reg_171][12  ( .D(D_12), .E(n6342), .C(wclk), .QN(n2028) );
  DFE1 \mem_reg_171][11  ( .D(D_11), .E(n6342), .C(wclk), .QN(n2029) );
  DFE1 \mem_reg_171][10  ( .D(D_10), .E(n6342), .C(wclk), .QN(n2030) );
  DFE1 \mem_reg_171][9  ( .D(D_9), .E(n6342), .C(wclk), .QN(n2031) );
  DFE1 \mem_reg_171][8  ( .D(D_8), .E(n6342), .C(wclk), .QN(n2032) );
  DFE1 \mem_reg_171][7  ( .D(D_7), .E(n6342), .C(wclk), .QN(n2033) );
  DFE1 \mem_reg_171][6  ( .D(D_6), .E(n6342), .C(wclk), .QN(n2034) );
  DFE1 \mem_reg_171][5  ( .D(D_5), .E(n6342), .C(wclk), .QN(n2035) );
  DFE1 \mem_reg_171][4  ( .D(D_4), .E(n6342), .C(wclk), .QN(n2036) );
  DFE1 \mem_reg_171][3  ( .D(D_3), .E(n6342), .C(wclk), .QN(n2037) );
  DFE1 \mem_reg_171][2  ( .D(D_2), .E(n6342), .C(wclk), .QN(n2038) );
  DFE1 \mem_reg_171][1  ( .D(D_1), .E(n6342), .C(wclk), .QN(n2039) );
  DFE1 \mem_reg_171][0  ( .D(D_0), .E(n6342), .C(wclk), .QN(n2040) );
  DFE1 \mem_reg_170][23  ( .D(D_23), .E(n6341), .C(wclk), .QN(n2041) );
  DFE1 \mem_reg_170][22  ( .D(D_22), .E(n6341), .C(wclk), .QN(n2042) );
  DFE1 \mem_reg_170][21  ( .D(D_21), .E(n6341), .C(wclk), .QN(n2043) );
  DFE1 \mem_reg_170][20  ( .D(D_20), .E(n6341), .C(wclk), .QN(n2044) );
  DFE1 \mem_reg_170][19  ( .D(D_19), .E(n6341), .C(wclk), .QN(n2045) );
  DFE1 \mem_reg_170][18  ( .D(D_18), .E(n6341), .C(wclk), .QN(n2046) );
  DFE1 \mem_reg_170][17  ( .D(D_17), .E(n6341), .C(wclk), .QN(n2047) );
  DFE1 \mem_reg_170][16  ( .D(D_16), .E(n6341), .C(wclk), .QN(n2048) );
  DFE1 \mem_reg_170][15  ( .D(D_15), .E(n6341), .C(wclk), .QN(n2049) );
  DFE1 \mem_reg_170][14  ( .D(D_14), .E(n6341), .C(wclk), .QN(n2050) );
  DFE1 \mem_reg_170][13  ( .D(D_13), .E(n6341), .C(wclk), .QN(n2051) );
  DFE1 \mem_reg_170][12  ( .D(D_12), .E(n6341), .C(wclk), .QN(n2052) );
  DFE1 \mem_reg_170][11  ( .D(D_11), .E(n6341), .C(wclk), .QN(n2053) );
  DFE1 \mem_reg_170][10  ( .D(D_10), .E(n6341), .C(wclk), .QN(n2054) );
  DFE1 \mem_reg_170][9  ( .D(D_9), .E(n6341), .C(wclk), .QN(n2055) );
  DFE1 \mem_reg_170][8  ( .D(D_8), .E(n6341), .C(wclk), .QN(n2056) );
  DFE1 \mem_reg_170][7  ( .D(D_7), .E(n6341), .C(wclk), .QN(n2057) );
  DFE1 \mem_reg_170][6  ( .D(D_6), .E(n6341), .C(wclk), .QN(n2058) );
  DFE1 \mem_reg_170][5  ( .D(D_5), .E(n6341), .C(wclk), .QN(n2059) );
  DFE1 \mem_reg_170][4  ( .D(D_4), .E(n6341), .C(wclk), .QN(n2060) );
  DFE1 \mem_reg_170][3  ( .D(D_3), .E(n6341), .C(wclk), .QN(n2061) );
  DFE1 \mem_reg_170][2  ( .D(D_2), .E(n6341), .C(wclk), .QN(n2062) );
  DFE1 \mem_reg_170][1  ( .D(D_1), .E(n6341), .C(wclk), .QN(n2063) );
  DFE1 \mem_reg_170][0  ( .D(D_0), .E(n6341), .C(wclk), .QN(n2064) );
  DFE1 \mem_reg_169][23  ( .D(D_23), .E(n6340), .C(wclk), .QN(n2065) );
  DFE1 \mem_reg_169][22  ( .D(D_22), .E(n6340), .C(wclk), .QN(n2066) );
  DFE1 \mem_reg_169][21  ( .D(D_21), .E(n6340), .C(wclk), .QN(n2067) );
  DFE1 \mem_reg_169][20  ( .D(D_20), .E(n6340), .C(wclk), .QN(n2068) );
  DFE1 \mem_reg_169][19  ( .D(D_19), .E(n6340), .C(wclk), .QN(n2069) );
  DFE1 \mem_reg_169][18  ( .D(D_18), .E(n6340), .C(wclk), .QN(n2070) );
  DFE1 \mem_reg_169][17  ( .D(D_17), .E(n6340), .C(wclk), .QN(n2071) );
  DFE1 \mem_reg_169][16  ( .D(D_16), .E(n6340), .C(wclk), .QN(n2072) );
  DFE1 \mem_reg_169][15  ( .D(D_15), .E(n6340), .C(wclk), .QN(n2073) );
  DFE1 \mem_reg_169][14  ( .D(D_14), .E(n6340), .C(wclk), .QN(n2074) );
  DFE1 \mem_reg_169][13  ( .D(D_13), .E(n6340), .C(wclk), .QN(n2075) );
  DFE1 \mem_reg_169][12  ( .D(D_12), .E(n6340), .C(wclk), .QN(n2076) );
  DFE1 \mem_reg_169][11  ( .D(D_11), .E(n6340), .C(wclk), .QN(n2077) );
  DFE1 \mem_reg_169][10  ( .D(D_10), .E(n6340), .C(wclk), .QN(n2078) );
  DFE1 \mem_reg_169][9  ( .D(D_9), .E(n6340), .C(wclk), .QN(n2079) );
  DFE1 \mem_reg_169][8  ( .D(D_8), .E(n6340), .C(wclk), .QN(n2080) );
  DFE1 \mem_reg_169][7  ( .D(D_7), .E(n6340), .C(wclk), .QN(n2081) );
  DFE1 \mem_reg_169][6  ( .D(D_6), .E(n6340), .C(wclk), .QN(n2082) );
  DFE1 \mem_reg_169][5  ( .D(D_5), .E(n6340), .C(wclk), .QN(n2083) );
  DFE1 \mem_reg_169][4  ( .D(D_4), .E(n6340), .C(wclk), .QN(n2084) );
  DFE1 \mem_reg_169][3  ( .D(D_3), .E(n6340), .C(wclk), .QN(n2085) );
  DFE1 \mem_reg_169][2  ( .D(D_2), .E(n6340), .C(wclk), .QN(n2086) );
  DFE1 \mem_reg_169][1  ( .D(D_1), .E(n6340), .C(wclk), .QN(n2087) );
  DFE1 \mem_reg_169][0  ( .D(D_0), .E(n6340), .C(wclk), .QN(n2088) );
  DFE1 \mem_reg_168][23  ( .D(D_23), .E(n6339), .C(wclk), .QN(n2089) );
  DFE1 \mem_reg_168][22  ( .D(D_22), .E(n6339), .C(wclk), .QN(n2090) );
  DFE1 \mem_reg_168][21  ( .D(D_21), .E(n6339), .C(wclk), .QN(n2091) );
  DFE1 \mem_reg_168][20  ( .D(D_20), .E(n6339), .C(wclk), .QN(n2092) );
  DFE1 \mem_reg_168][19  ( .D(D_19), .E(n6339), .C(wclk), .QN(n2093) );
  DFE1 \mem_reg_168][18  ( .D(D_18), .E(n6339), .C(wclk), .QN(n2094) );
  DFE1 \mem_reg_168][17  ( .D(D_17), .E(n6339), .C(wclk), .QN(n2095) );
  DFE1 \mem_reg_168][16  ( .D(D_16), .E(n6339), .C(wclk), .QN(n2096) );
  DFE1 \mem_reg_168][15  ( .D(D_15), .E(n6339), .C(wclk), .QN(n2097) );
  DFE1 \mem_reg_168][14  ( .D(D_14), .E(n6339), .C(wclk), .QN(n2098) );
  DFE1 \mem_reg_168][13  ( .D(D_13), .E(n6339), .C(wclk), .QN(n2099) );
  DFE1 \mem_reg_168][12  ( .D(D_12), .E(n6339), .C(wclk), .QN(n2100) );
  DFE1 \mem_reg_168][11  ( .D(D_11), .E(n6339), .C(wclk), .QN(n2101) );
  DFE1 \mem_reg_168][10  ( .D(D_10), .E(n6339), .C(wclk), .QN(n2102) );
  DFE1 \mem_reg_168][9  ( .D(D_9), .E(n6339), .C(wclk), .QN(n2103) );
  DFE1 \mem_reg_168][8  ( .D(D_8), .E(n6339), .C(wclk), .QN(n2104) );
  DFE1 \mem_reg_168][7  ( .D(D_7), .E(n6339), .C(wclk), .QN(n2105) );
  DFE1 \mem_reg_168][6  ( .D(D_6), .E(n6339), .C(wclk), .QN(n2106) );
  DFE1 \mem_reg_168][5  ( .D(D_5), .E(n6339), .C(wclk), .QN(n2107) );
  DFE1 \mem_reg_168][4  ( .D(D_4), .E(n6339), .C(wclk), .QN(n2108) );
  DFE1 \mem_reg_168][3  ( .D(D_3), .E(n6339), .C(wclk), .QN(n2109) );
  DFE1 \mem_reg_168][2  ( .D(D_2), .E(n6339), .C(wclk), .QN(n2110) );
  DFE1 \mem_reg_168][1  ( .D(D_1), .E(n6339), .C(wclk), .QN(n2111) );
  DFE1 \mem_reg_168][0  ( .D(D_0), .E(n6339), .C(wclk), .QN(n2112) );
  DFE1 \mem_reg_167][23  ( .D(D_23), .E(n6338), .C(wclk), .QN(n2113) );
  DFE1 \mem_reg_167][22  ( .D(D_22), .E(n6338), .C(wclk), .QN(n2114) );
  DFE1 \mem_reg_167][21  ( .D(D_21), .E(n6338), .C(wclk), .QN(n2115) );
  DFE1 \mem_reg_167][20  ( .D(D_20), .E(n6338), .C(wclk), .QN(n2116) );
  DFE1 \mem_reg_167][19  ( .D(D_19), .E(n6338), .C(wclk), .QN(n2117) );
  DFE1 \mem_reg_167][18  ( .D(D_18), .E(n6338), .C(wclk), .QN(n2118) );
  DFE1 \mem_reg_167][17  ( .D(D_17), .E(n6338), .C(wclk), .QN(n2119) );
  DFE1 \mem_reg_167][16  ( .D(D_16), .E(n6338), .C(wclk), .QN(n2120) );
  DFE1 \mem_reg_167][15  ( .D(D_15), .E(n6338), .C(wclk), .QN(n2121) );
  DFE1 \mem_reg_167][14  ( .D(D_14), .E(n6338), .C(wclk), .QN(n2122) );
  DFE1 \mem_reg_167][13  ( .D(D_13), .E(n6338), .C(wclk), .QN(n2123) );
  DFE1 \mem_reg_167][12  ( .D(D_12), .E(n6338), .C(wclk), .QN(n2124) );
  DFE1 \mem_reg_167][11  ( .D(D_11), .E(n6338), .C(wclk), .QN(n2125) );
  DFE1 \mem_reg_167][10  ( .D(D_10), .E(n6338), .C(wclk), .QN(n2126) );
  DFE1 \mem_reg_167][9  ( .D(D_9), .E(n6338), .C(wclk), .QN(n2127) );
  DFE1 \mem_reg_167][8  ( .D(D_8), .E(n6338), .C(wclk), .QN(n2128) );
  DFE1 \mem_reg_167][7  ( .D(D_7), .E(n6338), .C(wclk), .QN(n2129) );
  DFE1 \mem_reg_167][6  ( .D(D_6), .E(n6338), .C(wclk), .QN(n2130) );
  DFE1 \mem_reg_167][5  ( .D(D_5), .E(n6338), .C(wclk), .QN(n2131) );
  DFE1 \mem_reg_167][4  ( .D(D_4), .E(n6338), .C(wclk), .QN(n2132) );
  DFE1 \mem_reg_167][3  ( .D(D_3), .E(n6338), .C(wclk), .QN(n2133) );
  DFE1 \mem_reg_167][2  ( .D(D_2), .E(n6338), .C(wclk), .QN(n2134) );
  DFE1 \mem_reg_167][1  ( .D(D_1), .E(n6338), .C(wclk), .QN(n2135) );
  DFE1 \mem_reg_167][0  ( .D(D_0), .E(n6338), .C(wclk), .QN(n2136) );
  DFE1 \mem_reg_166][23  ( .D(D_23), .E(n6337), .C(wclk), .QN(n2137) );
  DFE1 \mem_reg_166][22  ( .D(D_22), .E(n6337), .C(wclk), .QN(n2138) );
  DFE1 \mem_reg_166][21  ( .D(D_21), .E(n6337), .C(wclk), .QN(n2139) );
  DFE1 \mem_reg_166][20  ( .D(D_20), .E(n6337), .C(wclk), .QN(n2140) );
  DFE1 \mem_reg_166][19  ( .D(D_19), .E(n6337), .C(wclk), .QN(n2141) );
  DFE1 \mem_reg_166][18  ( .D(D_18), .E(n6337), .C(wclk), .QN(n2142) );
  DFE1 \mem_reg_166][17  ( .D(D_17), .E(n6337), .C(wclk), .QN(n2143) );
  DFE1 \mem_reg_166][16  ( .D(D_16), .E(n6337), .C(wclk), .QN(n2144) );
  DFE1 \mem_reg_166][15  ( .D(D_15), .E(n6337), .C(wclk), .QN(n2145) );
  DFE1 \mem_reg_166][14  ( .D(D_14), .E(n6337), .C(wclk), .QN(n2146) );
  DFE1 \mem_reg_166][13  ( .D(D_13), .E(n6337), .C(wclk), .QN(n2147) );
  DFE1 \mem_reg_166][12  ( .D(D_12), .E(n6337), .C(wclk), .QN(n2148) );
  DFE1 \mem_reg_166][11  ( .D(D_11), .E(n6337), .C(wclk), .QN(n2149) );
  DFE1 \mem_reg_166][10  ( .D(D_10), .E(n6337), .C(wclk), .QN(n2150) );
  DFE1 \mem_reg_166][9  ( .D(D_9), .E(n6337), .C(wclk), .QN(n2151) );
  DFE1 \mem_reg_166][8  ( .D(D_8), .E(n6337), .C(wclk), .QN(n2152) );
  DFE1 \mem_reg_166][7  ( .D(D_7), .E(n6337), .C(wclk), .QN(n2153) );
  DFE1 \mem_reg_166][6  ( .D(D_6), .E(n6337), .C(wclk), .QN(n2154) );
  DFE1 \mem_reg_166][5  ( .D(D_5), .E(n6337), .C(wclk), .QN(n2155) );
  DFE1 \mem_reg_166][4  ( .D(D_4), .E(n6337), .C(wclk), .QN(n2156) );
  DFE1 \mem_reg_166][3  ( .D(D_3), .E(n6337), .C(wclk), .QN(n2157) );
  DFE1 \mem_reg_166][2  ( .D(D_2), .E(n6337), .C(wclk), .QN(n2158) );
  DFE1 \mem_reg_166][1  ( .D(D_1), .E(n6337), .C(wclk), .QN(n2159) );
  DFE1 \mem_reg_166][0  ( .D(D_0), .E(n6337), .C(wclk), .QN(n2160) );
  DFE1 \mem_reg_165][23  ( .D(D_23), .E(n6336), .C(wclk), .QN(n2161) );
  DFE1 \mem_reg_165][22  ( .D(D_22), .E(n6336), .C(wclk), .QN(n2162) );
  DFE1 \mem_reg_165][21  ( .D(D_21), .E(n6336), .C(wclk), .QN(n2163) );
  DFE1 \mem_reg_165][20  ( .D(D_20), .E(n6336), .C(wclk), .QN(n2164) );
  DFE1 \mem_reg_165][19  ( .D(D_19), .E(n6336), .C(wclk), .QN(n2165) );
  DFE1 \mem_reg_165][18  ( .D(D_18), .E(n6336), .C(wclk), .QN(n2166) );
  DFE1 \mem_reg_165][17  ( .D(D_17), .E(n6336), .C(wclk), .QN(n2167) );
  DFE1 \mem_reg_165][16  ( .D(D_16), .E(n6336), .C(wclk), .QN(n2168) );
  DFE1 \mem_reg_165][15  ( .D(D_15), .E(n6336), .C(wclk), .QN(n2169) );
  DFE1 \mem_reg_165][14  ( .D(D_14), .E(n6336), .C(wclk), .QN(n2170) );
  DFE1 \mem_reg_165][13  ( .D(D_13), .E(n6336), .C(wclk), .QN(n2171) );
  DFE1 \mem_reg_165][12  ( .D(D_12), .E(n6336), .C(wclk), .QN(n2172) );
  DFE1 \mem_reg_165][11  ( .D(D_11), .E(n6336), .C(wclk), .QN(n2173) );
  DFE1 \mem_reg_165][10  ( .D(D_10), .E(n6336), .C(wclk), .QN(n2174) );
  DFE1 \mem_reg_165][9  ( .D(D_9), .E(n6336), .C(wclk), .QN(n2175) );
  DFE1 \mem_reg_165][8  ( .D(D_8), .E(n6336), .C(wclk), .QN(n2176) );
  DFE1 \mem_reg_165][7  ( .D(D_7), .E(n6336), .C(wclk), .QN(n2177) );
  DFE1 \mem_reg_165][6  ( .D(D_6), .E(n6336), .C(wclk), .QN(n2178) );
  DFE1 \mem_reg_165][5  ( .D(D_5), .E(n6336), .C(wclk), .QN(n2179) );
  DFE1 \mem_reg_165][4  ( .D(D_4), .E(n6336), .C(wclk), .QN(n2180) );
  DFE1 \mem_reg_165][3  ( .D(D_3), .E(n6336), .C(wclk), .QN(n2181) );
  DFE1 \mem_reg_165][2  ( .D(D_2), .E(n6336), .C(wclk), .QN(n2182) );
  DFE1 \mem_reg_165][1  ( .D(D_1), .E(n6336), .C(wclk), .QN(n2183) );
  DFE1 \mem_reg_165][0  ( .D(D_0), .E(n6336), .C(wclk), .QN(n2184) );
  DFE1 \mem_reg_164][23  ( .D(D_23), .E(n6335), .C(wclk), .QN(n2185) );
  DFE1 \mem_reg_164][22  ( .D(D_22), .E(n6335), .C(wclk), .QN(n2186) );
  DFE1 \mem_reg_164][21  ( .D(D_21), .E(n6335), .C(wclk), .QN(n2187) );
  DFE1 \mem_reg_164][20  ( .D(D_20), .E(n6335), .C(wclk), .QN(n2188) );
  DFE1 \mem_reg_164][19  ( .D(D_19), .E(n6335), .C(wclk), .QN(n2189) );
  DFE1 \mem_reg_164][18  ( .D(D_18), .E(n6335), .C(wclk), .QN(n2190) );
  DFE1 \mem_reg_164][17  ( .D(D_17), .E(n6335), .C(wclk), .QN(n2191) );
  DFE1 \mem_reg_164][16  ( .D(D_16), .E(n6335), .C(wclk), .QN(n2192) );
  DFE1 \mem_reg_164][15  ( .D(D_15), .E(n6335), .C(wclk), .QN(n2193) );
  DFE1 \mem_reg_164][14  ( .D(D_14), .E(n6335), .C(wclk), .QN(n2194) );
  DFE1 \mem_reg_164][13  ( .D(D_13), .E(n6335), .C(wclk), .QN(n2195) );
  DFE1 \mem_reg_164][12  ( .D(D_12), .E(n6335), .C(wclk), .QN(n2196) );
  DFE1 \mem_reg_164][11  ( .D(D_11), .E(n6335), .C(wclk), .QN(n2197) );
  DFE1 \mem_reg_164][10  ( .D(D_10), .E(n6335), .C(wclk), .QN(n2198) );
  DFE1 \mem_reg_164][9  ( .D(D_9), .E(n6335), .C(wclk), .QN(n2199) );
  DFE1 \mem_reg_164][8  ( .D(D_8), .E(n6335), .C(wclk), .QN(n2200) );
  DFE1 \mem_reg_164][7  ( .D(D_7), .E(n6335), .C(wclk), .QN(n2201) );
  DFE1 \mem_reg_164][6  ( .D(D_6), .E(n6335), .C(wclk), .QN(n2202) );
  DFE1 \mem_reg_164][5  ( .D(D_5), .E(n6335), .C(wclk), .QN(n2203) );
  DFE1 \mem_reg_164][4  ( .D(D_4), .E(n6335), .C(wclk), .QN(n2204) );
  DFE1 \mem_reg_164][3  ( .D(D_3), .E(n6335), .C(wclk), .QN(n2205) );
  DFE1 \mem_reg_164][2  ( .D(D_2), .E(n6335), .C(wclk), .QN(n2206) );
  DFE1 \mem_reg_164][1  ( .D(D_1), .E(n6335), .C(wclk), .QN(n2207) );
  DFE1 \mem_reg_164][0  ( .D(D_0), .E(n6335), .C(wclk), .QN(n2208) );
  DFE1 \mem_reg_163][23  ( .D(D_23), .E(n6334), .C(wclk), .QN(n2209) );
  DFE1 \mem_reg_163][22  ( .D(D_22), .E(n6334), .C(wclk), .QN(n2210) );
  DFE1 \mem_reg_163][21  ( .D(D_21), .E(n6334), .C(wclk), .QN(n2211) );
  DFE1 \mem_reg_163][20  ( .D(D_20), .E(n6334), .C(wclk), .QN(n2212) );
  DFE1 \mem_reg_163][19  ( .D(D_19), .E(n6334), .C(wclk), .QN(n2213) );
  DFE1 \mem_reg_163][18  ( .D(D_18), .E(n6334), .C(wclk), .QN(n2214) );
  DFE1 \mem_reg_163][17  ( .D(D_17), .E(n6334), .C(wclk), .QN(n2215) );
  DFE1 \mem_reg_163][16  ( .D(D_16), .E(n6334), .C(wclk), .QN(n2216) );
  DFE1 \mem_reg_163][15  ( .D(D_15), .E(n6334), .C(wclk), .QN(n2217) );
  DFE1 \mem_reg_163][14  ( .D(D_14), .E(n6334), .C(wclk), .QN(n2218) );
  DFE1 \mem_reg_163][13  ( .D(D_13), .E(n6334), .C(wclk), .QN(n2219) );
  DFE1 \mem_reg_163][12  ( .D(D_12), .E(n6334), .C(wclk), .QN(n2220) );
  DFE1 \mem_reg_163][11  ( .D(D_11), .E(n6334), .C(wclk), .QN(n2221) );
  DFE1 \mem_reg_163][10  ( .D(D_10), .E(n6334), .C(wclk), .QN(n2222) );
  DFE1 \mem_reg_163][9  ( .D(D_9), .E(n6334), .C(wclk), .QN(n2223) );
  DFE1 \mem_reg_163][8  ( .D(D_8), .E(n6334), .C(wclk), .QN(n2224) );
  DFE1 \mem_reg_163][7  ( .D(D_7), .E(n6334), .C(wclk), .QN(n2225) );
  DFE1 \mem_reg_163][6  ( .D(D_6), .E(n6334), .C(wclk), .QN(n2226) );
  DFE1 \mem_reg_163][5  ( .D(D_5), .E(n6334), .C(wclk), .QN(n2227) );
  DFE1 \mem_reg_163][4  ( .D(D_4), .E(n6334), .C(wclk), .QN(n2228) );
  DFE1 \mem_reg_163][3  ( .D(D_3), .E(n6334), .C(wclk), .QN(n2229) );
  DFE1 \mem_reg_163][2  ( .D(D_2), .E(n6334), .C(wclk), .QN(n2230) );
  DFE1 \mem_reg_163][1  ( .D(D_1), .E(n6334), .C(wclk), .QN(n2231) );
  DFE1 \mem_reg_163][0  ( .D(D_0), .E(n6334), .C(wclk), .QN(n2232) );
  DFE1 \mem_reg_162][23  ( .D(D_23), .E(n6333), .C(wclk), .QN(n2233) );
  DFE1 \mem_reg_162][22  ( .D(D_22), .E(n6333), .C(wclk), .QN(n2234) );
  DFE1 \mem_reg_162][21  ( .D(D_21), .E(n6333), .C(wclk), .QN(n2235) );
  DFE1 \mem_reg_162][20  ( .D(D_20), .E(n6333), .C(wclk), .QN(n2236) );
  DFE1 \mem_reg_162][19  ( .D(D_19), .E(n6333), .C(wclk), .QN(n2237) );
  DFE1 \mem_reg_162][18  ( .D(D_18), .E(n6333), .C(wclk), .QN(n2238) );
  DFE1 \mem_reg_162][17  ( .D(D_17), .E(n6333), .C(wclk), .QN(n2239) );
  DFE1 \mem_reg_162][16  ( .D(D_16), .E(n6333), .C(wclk), .QN(n2240) );
  DFE1 \mem_reg_162][15  ( .D(D_15), .E(n6333), .C(wclk), .QN(n2241) );
  DFE1 \mem_reg_162][14  ( .D(D_14), .E(n6333), .C(wclk), .QN(n2242) );
  DFE1 \mem_reg_162][13  ( .D(D_13), .E(n6333), .C(wclk), .QN(n2243) );
  DFE1 \mem_reg_162][12  ( .D(D_12), .E(n6333), .C(wclk), .QN(n2244) );
  DFE1 \mem_reg_162][11  ( .D(D_11), .E(n6333), .C(wclk), .QN(n2245) );
  DFE1 \mem_reg_162][10  ( .D(D_10), .E(n6333), .C(wclk), .QN(n2246) );
  DFE1 \mem_reg_162][9  ( .D(D_9), .E(n6333), .C(wclk), .QN(n2247) );
  DFE1 \mem_reg_162][8  ( .D(D_8), .E(n6333), .C(wclk), .QN(n2248) );
  DFE1 \mem_reg_162][7  ( .D(D_7), .E(n6333), .C(wclk), .QN(n2249) );
  DFE1 \mem_reg_162][6  ( .D(D_6), .E(n6333), .C(wclk), .QN(n2250) );
  DFE1 \mem_reg_162][5  ( .D(D_5), .E(n6333), .C(wclk), .QN(n2251) );
  DFE1 \mem_reg_162][4  ( .D(D_4), .E(n6333), .C(wclk), .QN(n2252) );
  DFE1 \mem_reg_162][3  ( .D(D_3), .E(n6333), .C(wclk), .QN(n2253) );
  DFE1 \mem_reg_162][2  ( .D(D_2), .E(n6333), .C(wclk), .QN(n2254) );
  DFE1 \mem_reg_162][1  ( .D(D_1), .E(n6333), .C(wclk), .QN(n2255) );
  DFE1 \mem_reg_162][0  ( .D(D_0), .E(n6333), .C(wclk), .QN(n2256) );
  DFE1 \mem_reg_161][23  ( .D(D_23), .E(n6332), .C(wclk), .QN(n2257) );
  DFE1 \mem_reg_161][22  ( .D(D_22), .E(n6332), .C(wclk), .QN(n2258) );
  DFE1 \mem_reg_161][21  ( .D(D_21), .E(n6332), .C(wclk), .QN(n2259) );
  DFE1 \mem_reg_161][20  ( .D(D_20), .E(n6332), .C(wclk), .QN(n2260) );
  DFE1 \mem_reg_161][19  ( .D(D_19), .E(n6332), .C(wclk), .QN(n2261) );
  DFE1 \mem_reg_161][18  ( .D(D_18), .E(n6332), .C(wclk), .QN(n2262) );
  DFE1 \mem_reg_161][17  ( .D(D_17), .E(n6332), .C(wclk), .QN(n2263) );
  DFE1 \mem_reg_161][16  ( .D(D_16), .E(n6332), .C(wclk), .QN(n2264) );
  DFE1 \mem_reg_161][15  ( .D(D_15), .E(n6332), .C(wclk), .QN(n2265) );
  DFE1 \mem_reg_161][14  ( .D(D_14), .E(n6332), .C(wclk), .QN(n2266) );
  DFE1 \mem_reg_161][13  ( .D(D_13), .E(n6332), .C(wclk), .QN(n2267) );
  DFE1 \mem_reg_161][12  ( .D(D_12), .E(n6332), .C(wclk), .QN(n2268) );
  DFE1 \mem_reg_161][11  ( .D(D_11), .E(n6332), .C(wclk), .QN(n2269) );
  DFE1 \mem_reg_161][10  ( .D(D_10), .E(n6332), .C(wclk), .QN(n2270) );
  DFE1 \mem_reg_161][9  ( .D(D_9), .E(n6332), .C(wclk), .QN(n2271) );
  DFE1 \mem_reg_161][8  ( .D(D_8), .E(n6332), .C(wclk), .QN(n2272) );
  DFE1 \mem_reg_161][7  ( .D(D_7), .E(n6332), .C(wclk), .QN(n2273) );
  DFE1 \mem_reg_161][6  ( .D(D_6), .E(n6332), .C(wclk), .QN(n2274) );
  DFE1 \mem_reg_161][5  ( .D(D_5), .E(n6332), .C(wclk), .QN(n2275) );
  DFE1 \mem_reg_161][4  ( .D(D_4), .E(n6332), .C(wclk), .QN(n2276) );
  DFE1 \mem_reg_161][3  ( .D(D_3), .E(n6332), .C(wclk), .QN(n2277) );
  DFE1 \mem_reg_161][2  ( .D(D_2), .E(n6332), .C(wclk), .QN(n2278) );
  DFE1 \mem_reg_161][1  ( .D(D_1), .E(n6332), .C(wclk), .QN(n2279) );
  DFE1 \mem_reg_161][0  ( .D(D_0), .E(n6332), .C(wclk), .QN(n2280) );
  DFE1 \mem_reg_160][23  ( .D(D_23), .E(n6330), .C(wclk), .QN(n2281) );
  DFE1 \mem_reg_160][22  ( .D(D_22), .E(n6330), .C(wclk), .QN(n2282) );
  DFE1 \mem_reg_160][21  ( .D(D_21), .E(n6330), .C(wclk), .QN(n2283) );
  DFE1 \mem_reg_160][20  ( .D(D_20), .E(n6330), .C(wclk), .QN(n2284) );
  DFE1 \mem_reg_160][19  ( .D(D_19), .E(n6330), .C(wclk), .QN(n2285) );
  DFE1 \mem_reg_160][18  ( .D(D_18), .E(n6330), .C(wclk), .QN(n2286) );
  DFE1 \mem_reg_160][17  ( .D(D_17), .E(n6330), .C(wclk), .QN(n2287) );
  DFE1 \mem_reg_160][16  ( .D(D_16), .E(n6330), .C(wclk), .QN(n2288) );
  DFE1 \mem_reg_160][15  ( .D(D_15), .E(n6330), .C(wclk), .QN(n2289) );
  DFE1 \mem_reg_160][14  ( .D(D_14), .E(n6330), .C(wclk), .QN(n2290) );
  DFE1 \mem_reg_160][13  ( .D(D_13), .E(n6330), .C(wclk), .QN(n2291) );
  DFE1 \mem_reg_160][12  ( .D(D_12), .E(n6330), .C(wclk), .QN(n2292) );
  DFE1 \mem_reg_160][11  ( .D(D_11), .E(n6330), .C(wclk), .QN(n2293) );
  DFE1 \mem_reg_160][10  ( .D(D_10), .E(n6330), .C(wclk), .QN(n2294) );
  DFE1 \mem_reg_160][9  ( .D(D_9), .E(n6330), .C(wclk), .QN(n2295) );
  DFE1 \mem_reg_160][8  ( .D(D_8), .E(n6330), .C(wclk), .QN(n2296) );
  DFE1 \mem_reg_160][7  ( .D(D_7), .E(n6330), .C(wclk), .QN(n2297) );
  DFE1 \mem_reg_160][6  ( .D(D_6), .E(n6330), .C(wclk), .QN(n2298) );
  DFE1 \mem_reg_160][5  ( .D(D_5), .E(n6330), .C(wclk), .QN(n2299) );
  DFE1 \mem_reg_160][4  ( .D(D_4), .E(n6330), .C(wclk), .QN(n2300) );
  DFE1 \mem_reg_160][3  ( .D(D_3), .E(n6330), .C(wclk), .QN(n2301) );
  DFE1 \mem_reg_160][2  ( .D(D_2), .E(n6330), .C(wclk), .QN(n2302) );
  DFE1 \mem_reg_160][1  ( .D(D_1), .E(n6330), .C(wclk), .QN(n2303) );
  DFE1 \mem_reg_160][0  ( .D(D_0), .E(n6330), .C(wclk), .QN(n2304) );
  DFE1 \mem_reg_159][23  ( .D(D_23), .E(n6329), .C(wclk), .QN(n2305) );
  DFE1 \mem_reg_159][22  ( .D(D_22), .E(n6329), .C(wclk), .QN(n2306) );
  DFE1 \mem_reg_159][21  ( .D(D_21), .E(n6329), .C(wclk), .QN(n2307) );
  DFE1 \mem_reg_159][20  ( .D(D_20), .E(n6329), .C(wclk), .QN(n2308) );
  DFE1 \mem_reg_159][19  ( .D(D_19), .E(n6329), .C(wclk), .QN(n2309) );
  DFE1 \mem_reg_159][18  ( .D(D_18), .E(n6329), .C(wclk), .QN(n2310) );
  DFE1 \mem_reg_159][17  ( .D(D_17), .E(n6329), .C(wclk), .QN(n2311) );
  DFE1 \mem_reg_159][16  ( .D(D_16), .E(n6329), .C(wclk), .QN(n2312) );
  DFE1 \mem_reg_159][15  ( .D(D_15), .E(n6329), .C(wclk), .QN(n2313) );
  DFE1 \mem_reg_159][14  ( .D(D_14), .E(n6329), .C(wclk), .QN(n2314) );
  DFE1 \mem_reg_159][13  ( .D(D_13), .E(n6329), .C(wclk), .QN(n2315) );
  DFE1 \mem_reg_159][12  ( .D(D_12), .E(n6329), .C(wclk), .QN(n2316) );
  DFE1 \mem_reg_159][11  ( .D(D_11), .E(n6329), .C(wclk), .QN(n2317) );
  DFE1 \mem_reg_159][10  ( .D(D_10), .E(n6329), .C(wclk), .QN(n2318) );
  DFE1 \mem_reg_159][9  ( .D(D_9), .E(n6329), .C(wclk), .QN(n2319) );
  DFE1 \mem_reg_159][8  ( .D(D_8), .E(n6329), .C(wclk), .QN(n2320) );
  DFE1 \mem_reg_159][7  ( .D(D_7), .E(n6329), .C(wclk), .QN(n2321) );
  DFE1 \mem_reg_159][6  ( .D(D_6), .E(n6329), .C(wclk), .QN(n2322) );
  DFE1 \mem_reg_159][5  ( .D(D_5), .E(n6329), .C(wclk), .QN(n2323) );
  DFE1 \mem_reg_159][4  ( .D(D_4), .E(n6329), .C(wclk), .QN(n2324) );
  DFE1 \mem_reg_159][3  ( .D(D_3), .E(n6329), .C(wclk), .QN(n2325) );
  DFE1 \mem_reg_159][2  ( .D(D_2), .E(n6329), .C(wclk), .QN(n2326) );
  DFE1 \mem_reg_159][1  ( .D(D_1), .E(n6329), .C(wclk), .QN(n2327) );
  DFE1 \mem_reg_159][0  ( .D(D_0), .E(n6329), .C(wclk), .QN(n2328) );
  DFE1 \mem_reg_158][23  ( .D(D_23), .E(n6328), .C(wclk), .QN(n2329) );
  DFE1 \mem_reg_158][22  ( .D(D_22), .E(n6328), .C(wclk), .QN(n2330) );
  DFE1 \mem_reg_158][21  ( .D(D_21), .E(n6328), .C(wclk), .QN(n2331) );
  DFE1 \mem_reg_158][20  ( .D(D_20), .E(n6328), .C(wclk), .QN(n2332) );
  DFE1 \mem_reg_158][19  ( .D(D_19), .E(n6328), .C(wclk), .QN(n2333) );
  DFE1 \mem_reg_158][18  ( .D(D_18), .E(n6328), .C(wclk), .QN(n2334) );
  DFE1 \mem_reg_158][17  ( .D(D_17), .E(n6328), .C(wclk), .QN(n2335) );
  DFE1 \mem_reg_158][16  ( .D(D_16), .E(n6328), .C(wclk), .QN(n2336) );
  DFE1 \mem_reg_158][15  ( .D(D_15), .E(n6328), .C(wclk), .QN(n2337) );
  DFE1 \mem_reg_158][14  ( .D(D_14), .E(n6328), .C(wclk), .QN(n2338) );
  DFE1 \mem_reg_158][13  ( .D(D_13), .E(n6328), .C(wclk), .QN(n2339) );
  DFE1 \mem_reg_158][12  ( .D(D_12), .E(n6328), .C(wclk), .QN(n2340) );
  DFE1 \mem_reg_158][11  ( .D(D_11), .E(n6328), .C(wclk), .QN(n2341) );
  DFE1 \mem_reg_158][10  ( .D(D_10), .E(n6328), .C(wclk), .QN(n2342) );
  DFE1 \mem_reg_158][9  ( .D(D_9), .E(n6328), .C(wclk), .QN(n2343) );
  DFE1 \mem_reg_158][8  ( .D(D_8), .E(n6328), .C(wclk), .QN(n2344) );
  DFE1 \mem_reg_158][7  ( .D(D_7), .E(n6328), .C(wclk), .QN(n2345) );
  DFE1 \mem_reg_158][6  ( .D(D_6), .E(n6328), .C(wclk), .QN(n2346) );
  DFE1 \mem_reg_158][5  ( .D(D_5), .E(n6328), .C(wclk), .QN(n2347) );
  DFE1 \mem_reg_158][4  ( .D(D_4), .E(n6328), .C(wclk), .QN(n2348) );
  DFE1 \mem_reg_158][3  ( .D(D_3), .E(n6328), .C(wclk), .QN(n2349) );
  DFE1 \mem_reg_158][2  ( .D(D_2), .E(n6328), .C(wclk), .QN(n2350) );
  DFE1 \mem_reg_158][1  ( .D(D_1), .E(n6328), .C(wclk), .QN(n2351) );
  DFE1 \mem_reg_158][0  ( .D(D_0), .E(n6328), .C(wclk), .QN(n2352) );
  DFE1 \mem_reg_157][23  ( .D(D_23), .E(n6327), .C(wclk), .QN(n2353) );
  DFE1 \mem_reg_157][22  ( .D(D_22), .E(n6327), .C(wclk), .QN(n2354) );
  DFE1 \mem_reg_157][21  ( .D(D_21), .E(n6327), .C(wclk), .QN(n2355) );
  DFE1 \mem_reg_157][20  ( .D(D_20), .E(n6327), .C(wclk), .QN(n2356) );
  DFE1 \mem_reg_157][19  ( .D(D_19), .E(n6327), .C(wclk), .QN(n2357) );
  DFE1 \mem_reg_157][18  ( .D(D_18), .E(n6327), .C(wclk), .QN(n2358) );
  DFE1 \mem_reg_157][17  ( .D(D_17), .E(n6327), .C(wclk), .QN(n2359) );
  DFE1 \mem_reg_157][16  ( .D(D_16), .E(n6327), .C(wclk), .QN(n2360) );
  DFE1 \mem_reg_157][15  ( .D(D_15), .E(n6327), .C(wclk), .QN(n2361) );
  DFE1 \mem_reg_157][14  ( .D(D_14), .E(n6327), .C(wclk), .QN(n2362) );
  DFE1 \mem_reg_157][13  ( .D(D_13), .E(n6327), .C(wclk), .QN(n2363) );
  DFE1 \mem_reg_157][12  ( .D(D_12), .E(n6327), .C(wclk), .QN(n2364) );
  DFE1 \mem_reg_157][11  ( .D(D_11), .E(n6327), .C(wclk), .QN(n2365) );
  DFE1 \mem_reg_157][10  ( .D(D_10), .E(n6327), .C(wclk), .QN(n2366) );
  DFE1 \mem_reg_157][9  ( .D(D_9), .E(n6327), .C(wclk), .QN(n2367) );
  DFE1 \mem_reg_157][8  ( .D(D_8), .E(n6327), .C(wclk), .QN(n2368) );
  DFE1 \mem_reg_157][7  ( .D(D_7), .E(n6327), .C(wclk), .QN(n2369) );
  DFE1 \mem_reg_157][6  ( .D(D_6), .E(n6327), .C(wclk), .QN(n2370) );
  DFE1 \mem_reg_157][5  ( .D(D_5), .E(n6327), .C(wclk), .QN(n2371) );
  DFE1 \mem_reg_157][4  ( .D(D_4), .E(n6327), .C(wclk), .QN(n2372) );
  DFE1 \mem_reg_157][3  ( .D(D_3), .E(n6327), .C(wclk), .QN(n2373) );
  DFE1 \mem_reg_157][2  ( .D(D_2), .E(n6327), .C(wclk), .QN(n2374) );
  DFE1 \mem_reg_157][1  ( .D(D_1), .E(n6327), .C(wclk), .QN(n2375) );
  DFE1 \mem_reg_157][0  ( .D(D_0), .E(n6327), .C(wclk), .QN(n2376) );
  DFE1 \mem_reg_156][23  ( .D(D_23), .E(n6326), .C(wclk), .QN(n2377) );
  DFE1 \mem_reg_156][22  ( .D(D_22), .E(n6326), .C(wclk), .QN(n2378) );
  DFE1 \mem_reg_156][21  ( .D(D_21), .E(n6326), .C(wclk), .QN(n2379) );
  DFE1 \mem_reg_156][20  ( .D(D_20), .E(n6326), .C(wclk), .QN(n2380) );
  DFE1 \mem_reg_156][19  ( .D(D_19), .E(n6326), .C(wclk), .QN(n2381) );
  DFE1 \mem_reg_156][18  ( .D(D_18), .E(n6326), .C(wclk), .QN(n2382) );
  DFE1 \mem_reg_156][17  ( .D(D_17), .E(n6326), .C(wclk), .QN(n2383) );
  DFE1 \mem_reg_156][16  ( .D(D_16), .E(n6326), .C(wclk), .QN(n2384) );
  DFE1 \mem_reg_156][15  ( .D(D_15), .E(n6326), .C(wclk), .QN(n2385) );
  DFE1 \mem_reg_156][14  ( .D(D_14), .E(n6326), .C(wclk), .QN(n2386) );
  DFE1 \mem_reg_156][13  ( .D(D_13), .E(n6326), .C(wclk), .QN(n2387) );
  DFE1 \mem_reg_156][12  ( .D(D_12), .E(n6326), .C(wclk), .QN(n2388) );
  DFE1 \mem_reg_156][11  ( .D(D_11), .E(n6326), .C(wclk), .QN(n2389) );
  DFE1 \mem_reg_156][10  ( .D(D_10), .E(n6326), .C(wclk), .QN(n2390) );
  DFE1 \mem_reg_156][9  ( .D(D_9), .E(n6326), .C(wclk), .QN(n2391) );
  DFE1 \mem_reg_156][8  ( .D(D_8), .E(n6326), .C(wclk), .QN(n2392) );
  DFE1 \mem_reg_156][7  ( .D(D_7), .E(n6326), .C(wclk), .QN(n2393) );
  DFE1 \mem_reg_156][6  ( .D(D_6), .E(n6326), .C(wclk), .QN(n2394) );
  DFE1 \mem_reg_156][5  ( .D(D_5), .E(n6326), .C(wclk), .QN(n2395) );
  DFE1 \mem_reg_156][4  ( .D(D_4), .E(n6326), .C(wclk), .QN(n2396) );
  DFE1 \mem_reg_156][3  ( .D(D_3), .E(n6326), .C(wclk), .QN(n2397) );
  DFE1 \mem_reg_156][2  ( .D(D_2), .E(n6326), .C(wclk), .QN(n2398) );
  DFE1 \mem_reg_156][1  ( .D(D_1), .E(n6326), .C(wclk), .QN(n2399) );
  DFE1 \mem_reg_156][0  ( .D(D_0), .E(n6326), .C(wclk), .QN(n2400) );
  DFE1 \mem_reg_155][23  ( .D(D_23), .E(n6325), .C(wclk), .QN(n2401) );
  DFE1 \mem_reg_155][22  ( .D(D_22), .E(n6325), .C(wclk), .QN(n2402) );
  DFE1 \mem_reg_155][21  ( .D(D_21), .E(n6325), .C(wclk), .QN(n2403) );
  DFE1 \mem_reg_155][20  ( .D(D_20), .E(n6325), .C(wclk), .QN(n2404) );
  DFE1 \mem_reg_155][19  ( .D(D_19), .E(n6325), .C(wclk), .QN(n2405) );
  DFE1 \mem_reg_155][18  ( .D(D_18), .E(n6325), .C(wclk), .QN(n2406) );
  DFE1 \mem_reg_155][17  ( .D(D_17), .E(n6325), .C(wclk), .QN(n2407) );
  DFE1 \mem_reg_155][16  ( .D(D_16), .E(n6325), .C(wclk), .QN(n2408) );
  DFE1 \mem_reg_155][15  ( .D(D_15), .E(n6325), .C(wclk), .QN(n2409) );
  DFE1 \mem_reg_155][14  ( .D(D_14), .E(n6325), .C(wclk), .QN(n2410) );
  DFE1 \mem_reg_155][13  ( .D(D_13), .E(n6325), .C(wclk), .QN(n2411) );
  DFE1 \mem_reg_155][12  ( .D(D_12), .E(n6325), .C(wclk), .QN(n2412) );
  DFE1 \mem_reg_155][11  ( .D(D_11), .E(n6325), .C(wclk), .QN(n2413) );
  DFE1 \mem_reg_155][10  ( .D(D_10), .E(n6325), .C(wclk), .QN(n2414) );
  DFE1 \mem_reg_155][9  ( .D(D_9), .E(n6325), .C(wclk), .QN(n2415) );
  DFE1 \mem_reg_155][8  ( .D(D_8), .E(n6325), .C(wclk), .QN(n2416) );
  DFE1 \mem_reg_155][7  ( .D(D_7), .E(n6325), .C(wclk), .QN(n2417) );
  DFE1 \mem_reg_155][6  ( .D(D_6), .E(n6325), .C(wclk), .QN(n2418) );
  DFE1 \mem_reg_155][5  ( .D(D_5), .E(n6325), .C(wclk), .QN(n2419) );
  DFE1 \mem_reg_155][4  ( .D(D_4), .E(n6325), .C(wclk), .QN(n2420) );
  DFE1 \mem_reg_155][3  ( .D(D_3), .E(n6325), .C(wclk), .QN(n2421) );
  DFE1 \mem_reg_155][2  ( .D(D_2), .E(n6325), .C(wclk), .QN(n2422) );
  DFE1 \mem_reg_155][1  ( .D(D_1), .E(n6325), .C(wclk), .QN(n2423) );
  DFE1 \mem_reg_155][0  ( .D(D_0), .E(n6325), .C(wclk), .QN(n2424) );
  DFE1 \mem_reg_154][23  ( .D(D_23), .E(n6324), .C(wclk), .QN(n2425) );
  DFE1 \mem_reg_154][22  ( .D(D_22), .E(n6324), .C(wclk), .QN(n2426) );
  DFE1 \mem_reg_154][21  ( .D(D_21), .E(n6324), .C(wclk), .QN(n2427) );
  DFE1 \mem_reg_154][20  ( .D(D_20), .E(n6324), .C(wclk), .QN(n2428) );
  DFE1 \mem_reg_154][19  ( .D(D_19), .E(n6324), .C(wclk), .QN(n2429) );
  DFE1 \mem_reg_154][18  ( .D(D_18), .E(n6324), .C(wclk), .QN(n2430) );
  DFE1 \mem_reg_154][17  ( .D(D_17), .E(n6324), .C(wclk), .QN(n2431) );
  DFE1 \mem_reg_154][16  ( .D(D_16), .E(n6324), .C(wclk), .QN(n2432) );
  DFE1 \mem_reg_154][15  ( .D(D_15), .E(n6324), .C(wclk), .QN(n2433) );
  DFE1 \mem_reg_154][14  ( .D(D_14), .E(n6324), .C(wclk), .QN(n2434) );
  DFE1 \mem_reg_154][13  ( .D(D_13), .E(n6324), .C(wclk), .QN(n2435) );
  DFE1 \mem_reg_154][12  ( .D(D_12), .E(n6324), .C(wclk), .QN(n2436) );
  DFE1 \mem_reg_154][11  ( .D(D_11), .E(n6324), .C(wclk), .QN(n2437) );
  DFE1 \mem_reg_154][10  ( .D(D_10), .E(n6324), .C(wclk), .QN(n2438) );
  DFE1 \mem_reg_154][9  ( .D(D_9), .E(n6324), .C(wclk), .QN(n2439) );
  DFE1 \mem_reg_154][8  ( .D(D_8), .E(n6324), .C(wclk), .QN(n2440) );
  DFE1 \mem_reg_154][7  ( .D(D_7), .E(n6324), .C(wclk), .QN(n2441) );
  DFE1 \mem_reg_154][6  ( .D(D_6), .E(n6324), .C(wclk), .QN(n2442) );
  DFE1 \mem_reg_154][5  ( .D(D_5), .E(n6324), .C(wclk), .QN(n2443) );
  DFE1 \mem_reg_154][4  ( .D(D_4), .E(n6324), .C(wclk), .QN(n2444) );
  DFE1 \mem_reg_154][3  ( .D(D_3), .E(n6324), .C(wclk), .QN(n2445) );
  DFE1 \mem_reg_154][2  ( .D(D_2), .E(n6324), .C(wclk), .QN(n2446) );
  DFE1 \mem_reg_154][1  ( .D(D_1), .E(n6324), .C(wclk), .QN(n2447) );
  DFE1 \mem_reg_154][0  ( .D(D_0), .E(n6324), .C(wclk), .QN(n2448) );
  DFE1 \mem_reg_153][23  ( .D(D_23), .E(n6323), .C(wclk), .QN(n2449) );
  DFE1 \mem_reg_153][22  ( .D(D_22), .E(n6323), .C(wclk), .QN(n2450) );
  DFE1 \mem_reg_153][21  ( .D(D_21), .E(n6323), .C(wclk), .QN(n2451) );
  DFE1 \mem_reg_153][20  ( .D(D_20), .E(n6323), .C(wclk), .QN(n2452) );
  DFE1 \mem_reg_153][19  ( .D(D_19), .E(n6323), .C(wclk), .QN(n2453) );
  DFE1 \mem_reg_153][18  ( .D(D_18), .E(n6323), .C(wclk), .QN(n2454) );
  DFE1 \mem_reg_153][17  ( .D(D_17), .E(n6323), .C(wclk), .QN(n2455) );
  DFE1 \mem_reg_153][16  ( .D(D_16), .E(n6323), .C(wclk), .QN(n2456) );
  DFE1 \mem_reg_153][15  ( .D(D_15), .E(n6323), .C(wclk), .QN(n2457) );
  DFE1 \mem_reg_153][14  ( .D(D_14), .E(n6323), .C(wclk), .QN(n2458) );
  DFE1 \mem_reg_153][13  ( .D(D_13), .E(n6323), .C(wclk), .QN(n2459) );
  DFE1 \mem_reg_153][12  ( .D(D_12), .E(n6323), .C(wclk), .QN(n2460) );
  DFE1 \mem_reg_153][11  ( .D(D_11), .E(n6323), .C(wclk), .QN(n2461) );
  DFE1 \mem_reg_153][10  ( .D(D_10), .E(n6323), .C(wclk), .QN(n2462) );
  DFE1 \mem_reg_153][9  ( .D(D_9), .E(n6323), .C(wclk), .QN(n2463) );
  DFE1 \mem_reg_153][8  ( .D(D_8), .E(n6323), .C(wclk), .QN(n2464) );
  DFE1 \mem_reg_153][7  ( .D(D_7), .E(n6323), .C(wclk), .QN(n2465) );
  DFE1 \mem_reg_153][6  ( .D(D_6), .E(n6323), .C(wclk), .QN(n2466) );
  DFE1 \mem_reg_153][5  ( .D(D_5), .E(n6323), .C(wclk), .QN(n2467) );
  DFE1 \mem_reg_153][4  ( .D(D_4), .E(n6323), .C(wclk), .QN(n2468) );
  DFE1 \mem_reg_153][3  ( .D(D_3), .E(n6323), .C(wclk), .QN(n2469) );
  DFE1 \mem_reg_153][2  ( .D(D_2), .E(n6323), .C(wclk), .QN(n2470) );
  DFE1 \mem_reg_153][1  ( .D(D_1), .E(n6323), .C(wclk), .QN(n2471) );
  DFE1 \mem_reg_153][0  ( .D(D_0), .E(n6323), .C(wclk), .QN(n2472) );
  DFE1 \mem_reg_152][23  ( .D(D_23), .E(n6322), .C(wclk), .QN(n2473) );
  DFE1 \mem_reg_152][22  ( .D(D_22), .E(n6322), .C(wclk), .QN(n2474) );
  DFE1 \mem_reg_152][21  ( .D(D_21), .E(n6322), .C(wclk), .QN(n2475) );
  DFE1 \mem_reg_152][20  ( .D(D_20), .E(n6322), .C(wclk), .QN(n2476) );
  DFE1 \mem_reg_152][19  ( .D(D_19), .E(n6322), .C(wclk), .QN(n2477) );
  DFE1 \mem_reg_152][18  ( .D(D_18), .E(n6322), .C(wclk), .QN(n2478) );
  DFE1 \mem_reg_152][17  ( .D(D_17), .E(n6322), .C(wclk), .QN(n2479) );
  DFE1 \mem_reg_152][16  ( .D(D_16), .E(n6322), .C(wclk), .QN(n2480) );
  DFE1 \mem_reg_152][15  ( .D(D_15), .E(n6322), .C(wclk), .QN(n2481) );
  DFE1 \mem_reg_152][14  ( .D(D_14), .E(n6322), .C(wclk), .QN(n2482) );
  DFE1 \mem_reg_152][13  ( .D(D_13), .E(n6322), .C(wclk), .QN(n2483) );
  DFE1 \mem_reg_152][12  ( .D(D_12), .E(n6322), .C(wclk), .QN(n2484) );
  DFE1 \mem_reg_152][11  ( .D(D_11), .E(n6322), .C(wclk), .QN(n2485) );
  DFE1 \mem_reg_152][10  ( .D(D_10), .E(n6322), .C(wclk), .QN(n2486) );
  DFE1 \mem_reg_152][9  ( .D(D_9), .E(n6322), .C(wclk), .QN(n2487) );
  DFE1 \mem_reg_152][8  ( .D(D_8), .E(n6322), .C(wclk), .QN(n2488) );
  DFE1 \mem_reg_152][7  ( .D(D_7), .E(n6322), .C(wclk), .QN(n2489) );
  DFE1 \mem_reg_152][6  ( .D(D_6), .E(n6322), .C(wclk), .QN(n2490) );
  DFE1 \mem_reg_152][5  ( .D(D_5), .E(n6322), .C(wclk), .QN(n2491) );
  DFE1 \mem_reg_152][4  ( .D(D_4), .E(n6322), .C(wclk), .QN(n2492) );
  DFE1 \mem_reg_152][3  ( .D(D_3), .E(n6322), .C(wclk), .QN(n2493) );
  DFE1 \mem_reg_152][2  ( .D(D_2), .E(n6322), .C(wclk), .QN(n2494) );
  DFE1 \mem_reg_152][1  ( .D(D_1), .E(n6322), .C(wclk), .QN(n2495) );
  DFE1 \mem_reg_152][0  ( .D(D_0), .E(n6322), .C(wclk), .QN(n2496) );
  DFE1 \mem_reg_151][23  ( .D(D_23), .E(n6321), .C(wclk), .QN(n2497) );
  DFE1 \mem_reg_151][22  ( .D(D_22), .E(n6321), .C(wclk), .QN(n2498) );
  DFE1 \mem_reg_151][21  ( .D(D_21), .E(n6321), .C(wclk), .QN(n2499) );
  DFE1 \mem_reg_151][20  ( .D(D_20), .E(n6321), .C(wclk), .QN(n2500) );
  DFE1 \mem_reg_151][19  ( .D(D_19), .E(n6321), .C(wclk), .QN(n2501) );
  DFE1 \mem_reg_151][18  ( .D(D_18), .E(n6321), .C(wclk), .QN(n2502) );
  DFE1 \mem_reg_151][17  ( .D(D_17), .E(n6321), .C(wclk), .QN(n2503) );
  DFE1 \mem_reg_151][16  ( .D(D_16), .E(n6321), .C(wclk), .QN(n2504) );
  DFE1 \mem_reg_151][15  ( .D(D_15), .E(n6321), .C(wclk), .QN(n2505) );
  DFE1 \mem_reg_151][14  ( .D(D_14), .E(n6321), .C(wclk), .QN(n2506) );
  DFE1 \mem_reg_151][13  ( .D(D_13), .E(n6321), .C(wclk), .QN(n2507) );
  DFE1 \mem_reg_151][12  ( .D(D_12), .E(n6321), .C(wclk), .QN(n2508) );
  DFE1 \mem_reg_151][11  ( .D(D_11), .E(n6321), .C(wclk), .QN(n2509) );
  DFE1 \mem_reg_151][10  ( .D(D_10), .E(n6321), .C(wclk), .QN(n2510) );
  DFE1 \mem_reg_151][9  ( .D(D_9), .E(n6321), .C(wclk), .QN(n2511) );
  DFE1 \mem_reg_151][8  ( .D(D_8), .E(n6321), .C(wclk), .QN(n2512) );
  DFE1 \mem_reg_151][7  ( .D(D_7), .E(n6321), .C(wclk), .QN(n2513) );
  DFE1 \mem_reg_151][6  ( .D(D_6), .E(n6321), .C(wclk), .QN(n2514) );
  DFE1 \mem_reg_151][5  ( .D(D_5), .E(n6321), .C(wclk), .QN(n2515) );
  DFE1 \mem_reg_151][4  ( .D(D_4), .E(n6321), .C(wclk), .QN(n2516) );
  DFE1 \mem_reg_151][3  ( .D(D_3), .E(n6321), .C(wclk), .QN(n2517) );
  DFE1 \mem_reg_151][2  ( .D(D_2), .E(n6321), .C(wclk), .QN(n2518) );
  DFE1 \mem_reg_151][1  ( .D(D_1), .E(n6321), .C(wclk), .QN(n2519) );
  DFE1 \mem_reg_151][0  ( .D(D_0), .E(n6321), .C(wclk), .QN(n2520) );
  DFE1 \mem_reg_150][23  ( .D(D_23), .E(n6320), .C(wclk), .QN(n2521) );
  DFE1 \mem_reg_150][22  ( .D(D_22), .E(n6320), .C(wclk), .QN(n2522) );
  DFE1 \mem_reg_150][21  ( .D(D_21), .E(n6320), .C(wclk), .QN(n2523) );
  DFE1 \mem_reg_150][20  ( .D(D_20), .E(n6320), .C(wclk), .QN(n2524) );
  DFE1 \mem_reg_150][19  ( .D(D_19), .E(n6320), .C(wclk), .QN(n2525) );
  DFE1 \mem_reg_150][18  ( .D(D_18), .E(n6320), .C(wclk), .QN(n2526) );
  DFE1 \mem_reg_150][17  ( .D(D_17), .E(n6320), .C(wclk), .QN(n2527) );
  DFE1 \mem_reg_150][16  ( .D(D_16), .E(n6320), .C(wclk), .QN(n2528) );
  DFE1 \mem_reg_150][15  ( .D(D_15), .E(n6320), .C(wclk), .QN(n2529) );
  DFE1 \mem_reg_150][14  ( .D(D_14), .E(n6320), .C(wclk), .QN(n2530) );
  DFE1 \mem_reg_150][13  ( .D(D_13), .E(n6320), .C(wclk), .QN(n2531) );
  DFE1 \mem_reg_150][12  ( .D(D_12), .E(n6320), .C(wclk), .QN(n2532) );
  DFE1 \mem_reg_150][11  ( .D(D_11), .E(n6320), .C(wclk), .QN(n2533) );
  DFE1 \mem_reg_150][10  ( .D(D_10), .E(n6320), .C(wclk), .QN(n2534) );
  DFE1 \mem_reg_150][9  ( .D(D_9), .E(n6320), .C(wclk), .QN(n2535) );
  DFE1 \mem_reg_150][8  ( .D(D_8), .E(n6320), .C(wclk), .QN(n2536) );
  DFE1 \mem_reg_150][7  ( .D(D_7), .E(n6320), .C(wclk), .QN(n2537) );
  DFE1 \mem_reg_150][6  ( .D(D_6), .E(n6320), .C(wclk), .QN(n2538) );
  DFE1 \mem_reg_150][5  ( .D(D_5), .E(n6320), .C(wclk), .QN(n2539) );
  DFE1 \mem_reg_150][4  ( .D(D_4), .E(n6320), .C(wclk), .QN(n2540) );
  DFE1 \mem_reg_150][3  ( .D(D_3), .E(n6320), .C(wclk), .QN(n2541) );
  DFE1 \mem_reg_150][2  ( .D(D_2), .E(n6320), .C(wclk), .QN(n2542) );
  DFE1 \mem_reg_150][1  ( .D(D_1), .E(n6320), .C(wclk), .QN(n2543) );
  DFE1 \mem_reg_150][0  ( .D(D_0), .E(n6320), .C(wclk), .QN(n2544) );
  DFE1 \mem_reg_149][23  ( .D(D_23), .E(n6319), .C(wclk), .QN(n2545) );
  DFE1 \mem_reg_149][22  ( .D(D_22), .E(n6319), .C(wclk), .QN(n2546) );
  DFE1 \mem_reg_149][21  ( .D(D_21), .E(n6319), .C(wclk), .QN(n2547) );
  DFE1 \mem_reg_149][20  ( .D(D_20), .E(n6319), .C(wclk), .QN(n2548) );
  DFE1 \mem_reg_149][19  ( .D(D_19), .E(n6319), .C(wclk), .QN(n2549) );
  DFE1 \mem_reg_149][18  ( .D(D_18), .E(n6319), .C(wclk), .QN(n2550) );
  DFE1 \mem_reg_149][17  ( .D(D_17), .E(n6319), .C(wclk), .QN(n2551) );
  DFE1 \mem_reg_149][16  ( .D(D_16), .E(n6319), .C(wclk), .QN(n2552) );
  DFE1 \mem_reg_149][15  ( .D(D_15), .E(n6319), .C(wclk), .QN(n2553) );
  DFE1 \mem_reg_149][14  ( .D(D_14), .E(n6319), .C(wclk), .QN(n2554) );
  DFE1 \mem_reg_149][13  ( .D(D_13), .E(n6319), .C(wclk), .QN(n2555) );
  DFE1 \mem_reg_149][12  ( .D(D_12), .E(n6319), .C(wclk), .QN(n2556) );
  DFE1 \mem_reg_149][11  ( .D(D_11), .E(n6319), .C(wclk), .QN(n2557) );
  DFE1 \mem_reg_149][10  ( .D(D_10), .E(n6319), .C(wclk), .QN(n2558) );
  DFE1 \mem_reg_149][9  ( .D(D_9), .E(n6319), .C(wclk), .QN(n2559) );
  DFE1 \mem_reg_149][8  ( .D(D_8), .E(n6319), .C(wclk), .QN(n2560) );
  DFE1 \mem_reg_149][7  ( .D(D_7), .E(n6319), .C(wclk), .QN(n2561) );
  DFE1 \mem_reg_149][6  ( .D(D_6), .E(n6319), .C(wclk), .QN(n2562) );
  DFE1 \mem_reg_149][5  ( .D(D_5), .E(n6319), .C(wclk), .QN(n2563) );
  DFE1 \mem_reg_149][4  ( .D(D_4), .E(n6319), .C(wclk), .QN(n2564) );
  DFE1 \mem_reg_149][3  ( .D(D_3), .E(n6319), .C(wclk), .QN(n2565) );
  DFE1 \mem_reg_149][2  ( .D(D_2), .E(n6319), .C(wclk), .QN(n2566) );
  DFE1 \mem_reg_149][1  ( .D(D_1), .E(n6319), .C(wclk), .QN(n2567) );
  DFE1 \mem_reg_149][0  ( .D(D_0), .E(n6319), .C(wclk), .QN(n2568) );
  DFE1 \mem_reg_148][23  ( .D(D_23), .E(n6318), .C(wclk), .QN(n2569) );
  DFE1 \mem_reg_148][22  ( .D(D_22), .E(n6318), .C(wclk), .QN(n2570) );
  DFE1 \mem_reg_148][21  ( .D(D_21), .E(n6318), .C(wclk), .QN(n2571) );
  DFE1 \mem_reg_148][20  ( .D(D_20), .E(n6318), .C(wclk), .QN(n2572) );
  DFE1 \mem_reg_148][19  ( .D(D_19), .E(n6318), .C(wclk), .QN(n2573) );
  DFE1 \mem_reg_148][18  ( .D(D_18), .E(n6318), .C(wclk), .QN(n2574) );
  DFE1 \mem_reg_148][17  ( .D(D_17), .E(n6318), .C(wclk), .QN(n2575) );
  DFE1 \mem_reg_148][16  ( .D(D_16), .E(n6318), .C(wclk), .QN(n2576) );
  DFE1 \mem_reg_148][15  ( .D(D_15), .E(n6318), .C(wclk), .QN(n2577) );
  DFE1 \mem_reg_148][14  ( .D(D_14), .E(n6318), .C(wclk), .QN(n2578) );
  DFE1 \mem_reg_148][13  ( .D(D_13), .E(n6318), .C(wclk), .QN(n2579) );
  DFE1 \mem_reg_148][12  ( .D(D_12), .E(n6318), .C(wclk), .QN(n2580) );
  DFE1 \mem_reg_148][11  ( .D(D_11), .E(n6318), .C(wclk), .QN(n2581) );
  DFE1 \mem_reg_148][10  ( .D(D_10), .E(n6318), .C(wclk), .QN(n2582) );
  DFE1 \mem_reg_148][9  ( .D(D_9), .E(n6318), .C(wclk), .QN(n2583) );
  DFE1 \mem_reg_148][8  ( .D(D_8), .E(n6318), .C(wclk), .QN(n2584) );
  DFE1 \mem_reg_148][7  ( .D(D_7), .E(n6318), .C(wclk), .QN(n2585) );
  DFE1 \mem_reg_148][6  ( .D(D_6), .E(n6318), .C(wclk), .QN(n2586) );
  DFE1 \mem_reg_148][5  ( .D(D_5), .E(n6318), .C(wclk), .QN(n2587) );
  DFE1 \mem_reg_148][4  ( .D(D_4), .E(n6318), .C(wclk), .QN(n2588) );
  DFE1 \mem_reg_148][3  ( .D(D_3), .E(n6318), .C(wclk), .QN(n2589) );
  DFE1 \mem_reg_148][2  ( .D(D_2), .E(n6318), .C(wclk), .QN(n2590) );
  DFE1 \mem_reg_148][1  ( .D(D_1), .E(n6318), .C(wclk), .QN(n2591) );
  DFE1 \mem_reg_148][0  ( .D(D_0), .E(n6318), .C(wclk), .QN(n2592) );
  DFE1 \mem_reg_147][23  ( .D(D_23), .E(n6317), .C(wclk), .QN(n2593) );
  DFE1 \mem_reg_147][22  ( .D(D_22), .E(n6317), .C(wclk), .QN(n2594) );
  DFE1 \mem_reg_147][21  ( .D(D_21), .E(n6317), .C(wclk), .QN(n2595) );
  DFE1 \mem_reg_147][20  ( .D(D_20), .E(n6317), .C(wclk), .QN(n2596) );
  DFE1 \mem_reg_147][19  ( .D(D_19), .E(n6317), .C(wclk), .QN(n2597) );
  DFE1 \mem_reg_147][18  ( .D(D_18), .E(n6317), .C(wclk), .QN(n2598) );
  DFE1 \mem_reg_147][17  ( .D(D_17), .E(n6317), .C(wclk), .QN(n2599) );
  DFE1 \mem_reg_147][16  ( .D(D_16), .E(n6317), .C(wclk), .QN(n2600) );
  DFE1 \mem_reg_147][15  ( .D(D_15), .E(n6317), .C(wclk), .QN(n2601) );
  DFE1 \mem_reg_147][14  ( .D(D_14), .E(n6317), .C(wclk), .QN(n2602) );
  DFE1 \mem_reg_147][13  ( .D(D_13), .E(n6317), .C(wclk), .QN(n2603) );
  DFE1 \mem_reg_147][12  ( .D(D_12), .E(n6317), .C(wclk), .QN(n2604) );
  DFE1 \mem_reg_147][11  ( .D(D_11), .E(n6317), .C(wclk), .QN(n2605) );
  DFE1 \mem_reg_147][10  ( .D(D_10), .E(n6317), .C(wclk), .QN(n2606) );
  DFE1 \mem_reg_147][9  ( .D(D_9), .E(n6317), .C(wclk), .QN(n2607) );
  DFE1 \mem_reg_147][8  ( .D(D_8), .E(n6317), .C(wclk), .QN(n2608) );
  DFE1 \mem_reg_147][7  ( .D(D_7), .E(n6317), .C(wclk), .QN(n2609) );
  DFE1 \mem_reg_147][6  ( .D(D_6), .E(n6317), .C(wclk), .QN(n2610) );
  DFE1 \mem_reg_147][5  ( .D(D_5), .E(n6317), .C(wclk), .QN(n2611) );
  DFE1 \mem_reg_147][4  ( .D(D_4), .E(n6317), .C(wclk), .QN(n2612) );
  DFE1 \mem_reg_147][3  ( .D(D_3), .E(n6317), .C(wclk), .QN(n2613) );
  DFE1 \mem_reg_147][2  ( .D(D_2), .E(n6317), .C(wclk), .QN(n2614) );
  DFE1 \mem_reg_147][1  ( .D(D_1), .E(n6317), .C(wclk), .QN(n2615) );
  DFE1 \mem_reg_147][0  ( .D(D_0), .E(n6317), .C(wclk), .QN(n2616) );
  DFE1 \mem_reg_146][23  ( .D(D_23), .E(n6316), .C(wclk), .QN(n2617) );
  DFE1 \mem_reg_146][22  ( .D(D_22), .E(n6316), .C(wclk), .QN(n2618) );
  DFE1 \mem_reg_146][21  ( .D(D_21), .E(n6316), .C(wclk), .QN(n2619) );
  DFE1 \mem_reg_146][20  ( .D(D_20), .E(n6316), .C(wclk), .QN(n2620) );
  DFE1 \mem_reg_146][19  ( .D(D_19), .E(n6316), .C(wclk), .QN(n2621) );
  DFE1 \mem_reg_146][18  ( .D(D_18), .E(n6316), .C(wclk), .QN(n2622) );
  DFE1 \mem_reg_146][17  ( .D(D_17), .E(n6316), .C(wclk), .QN(n2623) );
  DFE1 \mem_reg_146][16  ( .D(D_16), .E(n6316), .C(wclk), .QN(n2624) );
  DFE1 \mem_reg_146][15  ( .D(D_15), .E(n6316), .C(wclk), .QN(n2625) );
  DFE1 \mem_reg_146][14  ( .D(D_14), .E(n6316), .C(wclk), .QN(n2626) );
  DFE1 \mem_reg_146][13  ( .D(D_13), .E(n6316), .C(wclk), .QN(n2627) );
  DFE1 \mem_reg_146][12  ( .D(D_12), .E(n6316), .C(wclk), .QN(n2628) );
  DFE1 \mem_reg_146][11  ( .D(D_11), .E(n6316), .C(wclk), .QN(n2629) );
  DFE1 \mem_reg_146][10  ( .D(D_10), .E(n6316), .C(wclk), .QN(n2630) );
  DFE1 \mem_reg_146][9  ( .D(D_9), .E(n6316), .C(wclk), .QN(n2631) );
  DFE1 \mem_reg_146][8  ( .D(D_8), .E(n6316), .C(wclk), .QN(n2632) );
  DFE1 \mem_reg_146][7  ( .D(D_7), .E(n6316), .C(wclk), .QN(n2633) );
  DFE1 \mem_reg_146][6  ( .D(D_6), .E(n6316), .C(wclk), .QN(n2634) );
  DFE1 \mem_reg_146][5  ( .D(D_5), .E(n6316), .C(wclk), .QN(n2635) );
  DFE1 \mem_reg_146][4  ( .D(D_4), .E(n6316), .C(wclk), .QN(n2636) );
  DFE1 \mem_reg_146][3  ( .D(D_3), .E(n6316), .C(wclk), .QN(n2637) );
  DFE1 \mem_reg_146][2  ( .D(D_2), .E(n6316), .C(wclk), .QN(n2638) );
  DFE1 \mem_reg_146][1  ( .D(D_1), .E(n6316), .C(wclk), .QN(n2639) );
  DFE1 \mem_reg_146][0  ( .D(D_0), .E(n6316), .C(wclk), .QN(n2640) );
  DFE1 \mem_reg_145][23  ( .D(D_23), .E(n6315), .C(wclk), .QN(n2641) );
  DFE1 \mem_reg_145][22  ( .D(D_22), .E(n6315), .C(wclk), .QN(n2642) );
  DFE1 \mem_reg_145][21  ( .D(D_21), .E(n6315), .C(wclk), .QN(n2643) );
  DFE1 \mem_reg_145][20  ( .D(D_20), .E(n6315), .C(wclk), .QN(n2644) );
  DFE1 \mem_reg_145][19  ( .D(D_19), .E(n6315), .C(wclk), .QN(n2645) );
  DFE1 \mem_reg_145][18  ( .D(D_18), .E(n6315), .C(wclk), .QN(n2646) );
  DFE1 \mem_reg_145][17  ( .D(D_17), .E(n6315), .C(wclk), .QN(n2647) );
  DFE1 \mem_reg_145][16  ( .D(D_16), .E(n6315), .C(wclk), .QN(n2648) );
  DFE1 \mem_reg_145][15  ( .D(D_15), .E(n6315), .C(wclk), .QN(n2649) );
  DFE1 \mem_reg_145][14  ( .D(D_14), .E(n6315), .C(wclk), .QN(n2650) );
  DFE1 \mem_reg_145][13  ( .D(D_13), .E(n6315), .C(wclk), .QN(n2651) );
  DFE1 \mem_reg_145][12  ( .D(D_12), .E(n6315), .C(wclk), .QN(n2652) );
  DFE1 \mem_reg_145][11  ( .D(D_11), .E(n6315), .C(wclk), .QN(n2653) );
  DFE1 \mem_reg_145][10  ( .D(D_10), .E(n6315), .C(wclk), .QN(n2654) );
  DFE1 \mem_reg_145][9  ( .D(D_9), .E(n6315), .C(wclk), .QN(n2655) );
  DFE1 \mem_reg_145][8  ( .D(D_8), .E(n6315), .C(wclk), .QN(n2656) );
  DFE1 \mem_reg_145][7  ( .D(D_7), .E(n6315), .C(wclk), .QN(n2657) );
  DFE1 \mem_reg_145][6  ( .D(D_6), .E(n6315), .C(wclk), .QN(n2658) );
  DFE1 \mem_reg_145][5  ( .D(D_5), .E(n6315), .C(wclk), .QN(n2659) );
  DFE1 \mem_reg_145][4  ( .D(D_4), .E(n6315), .C(wclk), .QN(n2660) );
  DFE1 \mem_reg_145][3  ( .D(D_3), .E(n6315), .C(wclk), .QN(n2661) );
  DFE1 \mem_reg_145][2  ( .D(D_2), .E(n6315), .C(wclk), .QN(n2662) );
  DFE1 \mem_reg_145][1  ( .D(D_1), .E(n6315), .C(wclk), .QN(n2663) );
  DFE1 \mem_reg_145][0  ( .D(D_0), .E(n6315), .C(wclk), .QN(n2664) );
  DFE1 \mem_reg_144][23  ( .D(D_23), .E(n6313), .C(wclk), .QN(n2665) );
  DFE1 \mem_reg_144][22  ( .D(D_22), .E(n6313), .C(wclk), .QN(n2666) );
  DFE1 \mem_reg_144][21  ( .D(D_21), .E(n6313), .C(wclk), .QN(n2667) );
  DFE1 \mem_reg_144][20  ( .D(D_20), .E(n6313), .C(wclk), .QN(n2668) );
  DFE1 \mem_reg_144][19  ( .D(D_19), .E(n6313), .C(wclk), .QN(n2669) );
  DFE1 \mem_reg_144][18  ( .D(D_18), .E(n6313), .C(wclk), .QN(n2670) );
  DFE1 \mem_reg_144][17  ( .D(D_17), .E(n6313), .C(wclk), .QN(n2671) );
  DFE1 \mem_reg_144][16  ( .D(D_16), .E(n6313), .C(wclk), .QN(n2672) );
  DFE1 \mem_reg_144][15  ( .D(D_15), .E(n6313), .C(wclk), .QN(n2673) );
  DFE1 \mem_reg_144][14  ( .D(D_14), .E(n6313), .C(wclk), .QN(n2674) );
  DFE1 \mem_reg_144][13  ( .D(D_13), .E(n6313), .C(wclk), .QN(n2675) );
  DFE1 \mem_reg_144][12  ( .D(D_12), .E(n6313), .C(wclk), .QN(n2676) );
  DFE1 \mem_reg_144][11  ( .D(D_11), .E(n6313), .C(wclk), .QN(n2677) );
  DFE1 \mem_reg_144][10  ( .D(D_10), .E(n6313), .C(wclk), .QN(n2678) );
  DFE1 \mem_reg_144][9  ( .D(D_9), .E(n6313), .C(wclk), .QN(n2679) );
  DFE1 \mem_reg_144][8  ( .D(D_8), .E(n6313), .C(wclk), .QN(n2680) );
  DFE1 \mem_reg_144][7  ( .D(D_7), .E(n6313), .C(wclk), .QN(n2681) );
  DFE1 \mem_reg_144][6  ( .D(D_6), .E(n6313), .C(wclk), .QN(n2682) );
  DFE1 \mem_reg_144][5  ( .D(D_5), .E(n6313), .C(wclk), .QN(n2683) );
  DFE1 \mem_reg_144][4  ( .D(D_4), .E(n6313), .C(wclk), .QN(n2684) );
  DFE1 \mem_reg_144][3  ( .D(D_3), .E(n6313), .C(wclk), .QN(n2685) );
  DFE1 \mem_reg_144][2  ( .D(D_2), .E(n6313), .C(wclk), .QN(n2686) );
  DFE1 \mem_reg_144][1  ( .D(D_1), .E(n6313), .C(wclk), .QN(n2687) );
  DFE1 \mem_reg_144][0  ( .D(D_0), .E(n6313), .C(wclk), .QN(n2688) );
  DFE1 \mem_reg_143][23  ( .D(D_23), .E(n6311), .C(wclk), .QN(n2689) );
  DFE1 \mem_reg_143][22  ( .D(D_22), .E(n6311), .C(wclk), .QN(n2690) );
  DFE1 \mem_reg_143][21  ( .D(D_21), .E(n6311), .C(wclk), .QN(n2691) );
  DFE1 \mem_reg_143][20  ( .D(D_20), .E(n6311), .C(wclk), .QN(n2692) );
  DFE1 \mem_reg_143][19  ( .D(D_19), .E(n6311), .C(wclk), .QN(n2693) );
  DFE1 \mem_reg_143][18  ( .D(D_18), .E(n6311), .C(wclk), .QN(n2694) );
  DFE1 \mem_reg_143][17  ( .D(D_17), .E(n6311), .C(wclk), .QN(n2695) );
  DFE1 \mem_reg_143][16  ( .D(D_16), .E(n6311), .C(wclk), .QN(n2696) );
  DFE1 \mem_reg_143][15  ( .D(D_15), .E(n6311), .C(wclk), .QN(n2697) );
  DFE1 \mem_reg_143][14  ( .D(D_14), .E(n6311), .C(wclk), .QN(n2698) );
  DFE1 \mem_reg_143][13  ( .D(D_13), .E(n6311), .C(wclk), .QN(n2699) );
  DFE1 \mem_reg_143][12  ( .D(D_12), .E(n6311), .C(wclk), .QN(n2700) );
  DFE1 \mem_reg_143][11  ( .D(D_11), .E(n6311), .C(wclk), .QN(n2701) );
  DFE1 \mem_reg_143][10  ( .D(D_10), .E(n6311), .C(wclk), .QN(n2702) );
  DFE1 \mem_reg_143][9  ( .D(D_9), .E(n6311), .C(wclk), .QN(n2703) );
  DFE1 \mem_reg_143][8  ( .D(D_8), .E(n6311), .C(wclk), .QN(n2704) );
  DFE1 \mem_reg_143][7  ( .D(D_7), .E(n6311), .C(wclk), .QN(n2705) );
  DFE1 \mem_reg_143][6  ( .D(D_6), .E(n6311), .C(wclk), .QN(n2706) );
  DFE1 \mem_reg_143][5  ( .D(D_5), .E(n6311), .C(wclk), .QN(n2707) );
  DFE1 \mem_reg_143][4  ( .D(D_4), .E(n6311), .C(wclk), .QN(n2708) );
  DFE1 \mem_reg_143][3  ( .D(D_3), .E(n6311), .C(wclk), .QN(n2709) );
  DFE1 \mem_reg_143][2  ( .D(D_2), .E(n6311), .C(wclk), .QN(n2710) );
  DFE1 \mem_reg_143][1  ( .D(D_1), .E(n6311), .C(wclk), .QN(n2711) );
  DFE1 \mem_reg_143][0  ( .D(D_0), .E(n6311), .C(wclk), .QN(n2712) );
  DFE1 \mem_reg_142][23  ( .D(D_23), .E(n6310), .C(wclk), .QN(n2713) );
  DFE1 \mem_reg_142][22  ( .D(D_22), .E(n6310), .C(wclk), .QN(n2714) );
  DFE1 \mem_reg_142][21  ( .D(D_21), .E(n6310), .C(wclk), .QN(n2715) );
  DFE1 \mem_reg_142][20  ( .D(D_20), .E(n6310), .C(wclk), .QN(n2716) );
  DFE1 \mem_reg_142][19  ( .D(D_19), .E(n6310), .C(wclk), .QN(n2717) );
  DFE1 \mem_reg_142][18  ( .D(D_18), .E(n6310), .C(wclk), .QN(n2718) );
  DFE1 \mem_reg_142][17  ( .D(D_17), .E(n6310), .C(wclk), .QN(n2719) );
  DFE1 \mem_reg_142][16  ( .D(D_16), .E(n6310), .C(wclk), .QN(n2720) );
  DFE1 \mem_reg_142][15  ( .D(D_15), .E(n6310), .C(wclk), .QN(n2721) );
  DFE1 \mem_reg_142][14  ( .D(D_14), .E(n6310), .C(wclk), .QN(n2722) );
  DFE1 \mem_reg_142][13  ( .D(D_13), .E(n6310), .C(wclk), .QN(n2723) );
  DFE1 \mem_reg_142][12  ( .D(D_12), .E(n6310), .C(wclk), .QN(n2724) );
  DFE1 \mem_reg_142][11  ( .D(D_11), .E(n6310), .C(wclk), .QN(n2725) );
  DFE1 \mem_reg_142][10  ( .D(D_10), .E(n6310), .C(wclk), .QN(n2726) );
  DFE1 \mem_reg_142][9  ( .D(D_9), .E(n6310), .C(wclk), .QN(n2727) );
  DFE1 \mem_reg_142][8  ( .D(D_8), .E(n6310), .C(wclk), .QN(n2728) );
  DFE1 \mem_reg_142][7  ( .D(D_7), .E(n6310), .C(wclk), .QN(n2729) );
  DFE1 \mem_reg_142][6  ( .D(D_6), .E(n6310), .C(wclk), .QN(n2730) );
  DFE1 \mem_reg_142][5  ( .D(D_5), .E(n6310), .C(wclk), .QN(n2731) );
  DFE1 \mem_reg_142][4  ( .D(D_4), .E(n6310), .C(wclk), .QN(n2732) );
  DFE1 \mem_reg_142][3  ( .D(D_3), .E(n6310), .C(wclk), .QN(n2733) );
  DFE1 \mem_reg_142][2  ( .D(D_2), .E(n6310), .C(wclk), .QN(n2734) );
  DFE1 \mem_reg_142][1  ( .D(D_1), .E(n6310), .C(wclk), .QN(n2735) );
  DFE1 \mem_reg_142][0  ( .D(D_0), .E(n6310), .C(wclk), .QN(n2736) );
  DFE1 \mem_reg_141][23  ( .D(D_23), .E(n6309), .C(wclk), .QN(n2737) );
  DFE1 \mem_reg_141][22  ( .D(D_22), .E(n6309), .C(wclk), .QN(n2738) );
  DFE1 \mem_reg_141][21  ( .D(D_21), .E(n6309), .C(wclk), .QN(n2739) );
  DFE1 \mem_reg_141][20  ( .D(D_20), .E(n6309), .C(wclk), .QN(n2740) );
  DFE1 \mem_reg_141][19  ( .D(D_19), .E(n6309), .C(wclk), .QN(n2741) );
  DFE1 \mem_reg_141][18  ( .D(D_18), .E(n6309), .C(wclk), .QN(n2742) );
  DFE1 \mem_reg_141][17  ( .D(D_17), .E(n6309), .C(wclk), .QN(n2743) );
  DFE1 \mem_reg_141][16  ( .D(D_16), .E(n6309), .C(wclk), .QN(n2744) );
  DFE1 \mem_reg_141][15  ( .D(D_15), .E(n6309), .C(wclk), .QN(n2745) );
  DFE1 \mem_reg_141][14  ( .D(D_14), .E(n6309), .C(wclk), .QN(n2746) );
  DFE1 \mem_reg_141][13  ( .D(D_13), .E(n6309), .C(wclk), .QN(n2747) );
  DFE1 \mem_reg_141][12  ( .D(D_12), .E(n6309), .C(wclk), .QN(n2748) );
  DFE1 \mem_reg_141][11  ( .D(D_11), .E(n6309), .C(wclk), .QN(n2749) );
  DFE1 \mem_reg_141][10  ( .D(D_10), .E(n6309), .C(wclk), .QN(n2750) );
  DFE1 \mem_reg_141][9  ( .D(D_9), .E(n6309), .C(wclk), .QN(n2751) );
  DFE1 \mem_reg_141][8  ( .D(D_8), .E(n6309), .C(wclk), .QN(n2752) );
  DFE1 \mem_reg_141][7  ( .D(D_7), .E(n6309), .C(wclk), .QN(n2753) );
  DFE1 \mem_reg_141][6  ( .D(D_6), .E(n6309), .C(wclk), .QN(n2754) );
  DFE1 \mem_reg_141][5  ( .D(D_5), .E(n6309), .C(wclk), .QN(n2755) );
  DFE1 \mem_reg_141][4  ( .D(D_4), .E(n6309), .C(wclk), .QN(n2756) );
  DFE1 \mem_reg_141][3  ( .D(D_3), .E(n6309), .C(wclk), .QN(n2757) );
  DFE1 \mem_reg_141][2  ( .D(D_2), .E(n6309), .C(wclk), .QN(n2758) );
  DFE1 \mem_reg_141][1  ( .D(D_1), .E(n6309), .C(wclk), .QN(n2759) );
  DFE1 \mem_reg_141][0  ( .D(D_0), .E(n6309), .C(wclk), .QN(n2760) );
  DFE1 \mem_reg_140][23  ( .D(D_23), .E(n6308), .C(wclk), .QN(n2761) );
  DFE1 \mem_reg_140][22  ( .D(D_22), .E(n6308), .C(wclk), .QN(n2762) );
  DFE1 \mem_reg_140][21  ( .D(D_21), .E(n6308), .C(wclk), .QN(n2763) );
  DFE1 \mem_reg_140][20  ( .D(D_20), .E(n6308), .C(wclk), .QN(n2764) );
  DFE1 \mem_reg_140][19  ( .D(D_19), .E(n6308), .C(wclk), .QN(n2765) );
  DFE1 \mem_reg_140][18  ( .D(D_18), .E(n6308), .C(wclk), .QN(n2766) );
  DFE1 \mem_reg_140][17  ( .D(D_17), .E(n6308), .C(wclk), .QN(n2767) );
  DFE1 \mem_reg_140][16  ( .D(D_16), .E(n6308), .C(wclk), .QN(n2768) );
  DFE1 \mem_reg_140][15  ( .D(D_15), .E(n6308), .C(wclk), .QN(n2769) );
  DFE1 \mem_reg_140][14  ( .D(D_14), .E(n6308), .C(wclk), .QN(n2770) );
  DFE1 \mem_reg_140][13  ( .D(D_13), .E(n6308), .C(wclk), .QN(n2771) );
  DFE1 \mem_reg_140][12  ( .D(D_12), .E(n6308), .C(wclk), .QN(n2772) );
  DFE1 \mem_reg_140][11  ( .D(D_11), .E(n6308), .C(wclk), .QN(n2773) );
  DFE1 \mem_reg_140][10  ( .D(D_10), .E(n6308), .C(wclk), .QN(n2774) );
  DFE1 \mem_reg_140][9  ( .D(D_9), .E(n6308), .C(wclk), .QN(n2775) );
  DFE1 \mem_reg_140][8  ( .D(D_8), .E(n6308), .C(wclk), .QN(n2776) );
  DFE1 \mem_reg_140][7  ( .D(D_7), .E(n6308), .C(wclk), .QN(n2777) );
  DFE1 \mem_reg_140][6  ( .D(D_6), .E(n6308), .C(wclk), .QN(n2778) );
  DFE1 \mem_reg_140][5  ( .D(D_5), .E(n6308), .C(wclk), .QN(n2779) );
  DFE1 \mem_reg_140][4  ( .D(D_4), .E(n6308), .C(wclk), .QN(n2780) );
  DFE1 \mem_reg_140][3  ( .D(D_3), .E(n6308), .C(wclk), .QN(n2781) );
  DFE1 \mem_reg_140][2  ( .D(D_2), .E(n6308), .C(wclk), .QN(n2782) );
  DFE1 \mem_reg_140][1  ( .D(D_1), .E(n6308), .C(wclk), .QN(n2783) );
  DFE1 \mem_reg_140][0  ( .D(D_0), .E(n6308), .C(wclk), .QN(n2784) );
  DFE1 \mem_reg_139][23  ( .D(D_23), .E(n6307), .C(wclk), .QN(n2785) );
  DFE1 \mem_reg_139][22  ( .D(D_22), .E(n6307), .C(wclk), .QN(n2786) );
  DFE1 \mem_reg_139][21  ( .D(D_21), .E(n6307), .C(wclk), .QN(n2787) );
  DFE1 \mem_reg_139][20  ( .D(D_20), .E(n6307), .C(wclk), .QN(n2788) );
  DFE1 \mem_reg_139][19  ( .D(D_19), .E(n6307), .C(wclk), .QN(n2789) );
  DFE1 \mem_reg_139][18  ( .D(D_18), .E(n6307), .C(wclk), .QN(n2790) );
  DFE1 \mem_reg_139][17  ( .D(D_17), .E(n6307), .C(wclk), .QN(n2791) );
  DFE1 \mem_reg_139][16  ( .D(D_16), .E(n6307), .C(wclk), .QN(n2792) );
  DFE1 \mem_reg_139][15  ( .D(D_15), .E(n6307), .C(wclk), .QN(n2793) );
  DFE1 \mem_reg_139][14  ( .D(D_14), .E(n6307), .C(wclk), .QN(n2794) );
  DFE1 \mem_reg_139][13  ( .D(D_13), .E(n6307), .C(wclk), .QN(n2795) );
  DFE1 \mem_reg_139][12  ( .D(D_12), .E(n6307), .C(wclk), .QN(n2796) );
  DFE1 \mem_reg_139][11  ( .D(D_11), .E(n6307), .C(wclk), .QN(n2797) );
  DFE1 \mem_reg_139][10  ( .D(D_10), .E(n6307), .C(wclk), .QN(n2798) );
  DFE1 \mem_reg_139][9  ( .D(D_9), .E(n6307), .C(wclk), .QN(n2799) );
  DFE1 \mem_reg_139][8  ( .D(D_8), .E(n6307), .C(wclk), .QN(n2800) );
  DFE1 \mem_reg_139][7  ( .D(D_7), .E(n6307), .C(wclk), .QN(n2801) );
  DFE1 \mem_reg_139][6  ( .D(D_6), .E(n6307), .C(wclk), .QN(n2802) );
  DFE1 \mem_reg_139][5  ( .D(D_5), .E(n6307), .C(wclk), .QN(n2803) );
  DFE1 \mem_reg_139][4  ( .D(D_4), .E(n6307), .C(wclk), .QN(n2804) );
  DFE1 \mem_reg_139][3  ( .D(D_3), .E(n6307), .C(wclk), .QN(n2805) );
  DFE1 \mem_reg_139][2  ( .D(D_2), .E(n6307), .C(wclk), .QN(n2806) );
  DFE1 \mem_reg_139][1  ( .D(D_1), .E(n6307), .C(wclk), .QN(n2807) );
  DFE1 \mem_reg_139][0  ( .D(D_0), .E(n6307), .C(wclk), .QN(n2808) );
  DFE1 \mem_reg_138][23  ( .D(D_23), .E(n6306), .C(wclk), .QN(n2809) );
  DFE1 \mem_reg_138][22  ( .D(D_22), .E(n6306), .C(wclk), .QN(n2810) );
  DFE1 \mem_reg_138][21  ( .D(D_21), .E(n6306), .C(wclk), .QN(n2811) );
  DFE1 \mem_reg_138][20  ( .D(D_20), .E(n6306), .C(wclk), .QN(n2812) );
  DFE1 \mem_reg_138][19  ( .D(D_19), .E(n6306), .C(wclk), .QN(n2813) );
  DFE1 \mem_reg_138][18  ( .D(D_18), .E(n6306), .C(wclk), .QN(n2814) );
  DFE1 \mem_reg_138][17  ( .D(D_17), .E(n6306), .C(wclk), .QN(n2815) );
  DFE1 \mem_reg_138][16  ( .D(D_16), .E(n6306), .C(wclk), .QN(n2816) );
  DFE1 \mem_reg_138][15  ( .D(D_15), .E(n6306), .C(wclk), .QN(n2817) );
  DFE1 \mem_reg_138][14  ( .D(D_14), .E(n6306), .C(wclk), .QN(n2818) );
  DFE1 \mem_reg_138][13  ( .D(D_13), .E(n6306), .C(wclk), .QN(n2819) );
  DFE1 \mem_reg_138][12  ( .D(D_12), .E(n6306), .C(wclk), .QN(n2820) );
  DFE1 \mem_reg_138][11  ( .D(D_11), .E(n6306), .C(wclk), .QN(n2821) );
  DFE1 \mem_reg_138][10  ( .D(D_10), .E(n6306), .C(wclk), .QN(n2822) );
  DFE1 \mem_reg_138][9  ( .D(D_9), .E(n6306), .C(wclk), .QN(n2823) );
  DFE1 \mem_reg_138][8  ( .D(D_8), .E(n6306), .C(wclk), .QN(n2824) );
  DFE1 \mem_reg_138][7  ( .D(D_7), .E(n6306), .C(wclk), .QN(n2825) );
  DFE1 \mem_reg_138][6  ( .D(D_6), .E(n6306), .C(wclk), .QN(n2826) );
  DFE1 \mem_reg_138][5  ( .D(D_5), .E(n6306), .C(wclk), .QN(n2827) );
  DFE1 \mem_reg_138][4  ( .D(D_4), .E(n6306), .C(wclk), .QN(n2828) );
  DFE1 \mem_reg_138][3  ( .D(D_3), .E(n6306), .C(wclk), .QN(n2829) );
  DFE1 \mem_reg_138][2  ( .D(D_2), .E(n6306), .C(wclk), .QN(n2830) );
  DFE1 \mem_reg_138][1  ( .D(D_1), .E(n6306), .C(wclk), .QN(n2831) );
  DFE1 \mem_reg_138][0  ( .D(D_0), .E(n6306), .C(wclk), .QN(n2832) );
  DFE1 \mem_reg_137][23  ( .D(D_23), .E(n6305), .C(wclk), .QN(n2833) );
  DFE1 \mem_reg_137][22  ( .D(D_22), .E(n6305), .C(wclk), .QN(n2834) );
  DFE1 \mem_reg_137][21  ( .D(D_21), .E(n6305), .C(wclk), .QN(n2835) );
  DFE1 \mem_reg_137][20  ( .D(D_20), .E(n6305), .C(wclk), .QN(n2836) );
  DFE1 \mem_reg_137][19  ( .D(D_19), .E(n6305), .C(wclk), .QN(n2837) );
  DFE1 \mem_reg_137][18  ( .D(D_18), .E(n6305), .C(wclk), .QN(n2838) );
  DFE1 \mem_reg_137][17  ( .D(D_17), .E(n6305), .C(wclk), .QN(n2839) );
  DFE1 \mem_reg_137][16  ( .D(D_16), .E(n6305), .C(wclk), .QN(n2840) );
  DFE1 \mem_reg_137][15  ( .D(D_15), .E(n6305), .C(wclk), .QN(n2841) );
  DFE1 \mem_reg_137][14  ( .D(D_14), .E(n6305), .C(wclk), .QN(n2842) );
  DFE1 \mem_reg_137][13  ( .D(D_13), .E(n6305), .C(wclk), .QN(n2843) );
  DFE1 \mem_reg_137][12  ( .D(D_12), .E(n6305), .C(wclk), .QN(n2844) );
  DFE1 \mem_reg_137][11  ( .D(D_11), .E(n6305), .C(wclk), .QN(n2845) );
  DFE1 \mem_reg_137][10  ( .D(D_10), .E(n6305), .C(wclk), .QN(n2846) );
  DFE1 \mem_reg_137][9  ( .D(D_9), .E(n6305), .C(wclk), .QN(n2847) );
  DFE1 \mem_reg_137][8  ( .D(D_8), .E(n6305), .C(wclk), .QN(n2848) );
  DFE1 \mem_reg_137][7  ( .D(D_7), .E(n6305), .C(wclk), .QN(n2849) );
  DFE1 \mem_reg_137][6  ( .D(D_6), .E(n6305), .C(wclk), .QN(n2850) );
  DFE1 \mem_reg_137][5  ( .D(D_5), .E(n6305), .C(wclk), .QN(n2851) );
  DFE1 \mem_reg_137][4  ( .D(D_4), .E(n6305), .C(wclk), .QN(n2852) );
  DFE1 \mem_reg_137][3  ( .D(D_3), .E(n6305), .C(wclk), .QN(n2853) );
  DFE1 \mem_reg_137][2  ( .D(D_2), .E(n6305), .C(wclk), .QN(n2854) );
  DFE1 \mem_reg_137][1  ( .D(D_1), .E(n6305), .C(wclk), .QN(n2855) );
  DFE1 \mem_reg_137][0  ( .D(D_0), .E(n6305), .C(wclk), .QN(n2856) );
  DFE1 \mem_reg_136][23  ( .D(D_23), .E(n6304), .C(wclk), .QN(n2857) );
  DFE1 \mem_reg_136][22  ( .D(D_22), .E(n6304), .C(wclk), .QN(n2858) );
  DFE1 \mem_reg_136][21  ( .D(D_21), .E(n6304), .C(wclk), .QN(n2859) );
  DFE1 \mem_reg_136][20  ( .D(D_20), .E(n6304), .C(wclk), .QN(n2860) );
  DFE1 \mem_reg_136][19  ( .D(D_19), .E(n6304), .C(wclk), .QN(n2861) );
  DFE1 \mem_reg_136][18  ( .D(D_18), .E(n6304), .C(wclk), .QN(n2862) );
  DFE1 \mem_reg_136][17  ( .D(D_17), .E(n6304), .C(wclk), .QN(n2863) );
  DFE1 \mem_reg_136][16  ( .D(D_16), .E(n6304), .C(wclk), .QN(n2864) );
  DFE1 \mem_reg_136][15  ( .D(D_15), .E(n6304), .C(wclk), .QN(n2865) );
  DFE1 \mem_reg_136][14  ( .D(D_14), .E(n6304), .C(wclk), .QN(n2866) );
  DFE1 \mem_reg_136][13  ( .D(D_13), .E(n6304), .C(wclk), .QN(n2867) );
  DFE1 \mem_reg_136][12  ( .D(D_12), .E(n6304), .C(wclk), .QN(n2868) );
  DFE1 \mem_reg_136][11  ( .D(D_11), .E(n6304), .C(wclk), .QN(n2869) );
  DFE1 \mem_reg_136][10  ( .D(D_10), .E(n6304), .C(wclk), .QN(n2870) );
  DFE1 \mem_reg_136][9  ( .D(D_9), .E(n6304), .C(wclk), .QN(n2871) );
  DFE1 \mem_reg_136][8  ( .D(D_8), .E(n6304), .C(wclk), .QN(n2872) );
  DFE1 \mem_reg_136][7  ( .D(D_7), .E(n6304), .C(wclk), .QN(n2873) );
  DFE1 \mem_reg_136][6  ( .D(D_6), .E(n6304), .C(wclk), .QN(n2874) );
  DFE1 \mem_reg_136][5  ( .D(D_5), .E(n6304), .C(wclk), .QN(n2875) );
  DFE1 \mem_reg_136][4  ( .D(D_4), .E(n6304), .C(wclk), .QN(n2876) );
  DFE1 \mem_reg_136][3  ( .D(D_3), .E(n6304), .C(wclk), .QN(n2877) );
  DFE1 \mem_reg_136][2  ( .D(D_2), .E(n6304), .C(wclk), .QN(n2878) );
  DFE1 \mem_reg_136][1  ( .D(D_1), .E(n6304), .C(wclk), .QN(n2879) );
  DFE1 \mem_reg_136][0  ( .D(D_0), .E(n6304), .C(wclk), .QN(n2880) );
  DFE1 \mem_reg_135][23  ( .D(D_23), .E(n6303), .C(wclk), .QN(n2881) );
  DFE1 \mem_reg_135][22  ( .D(D_22), .E(n6303), .C(wclk), .QN(n2882) );
  DFE1 \mem_reg_135][21  ( .D(D_21), .E(n6303), .C(wclk), .QN(n2883) );
  DFE1 \mem_reg_135][20  ( .D(D_20), .E(n6303), .C(wclk), .QN(n2884) );
  DFE1 \mem_reg_135][19  ( .D(D_19), .E(n6303), .C(wclk), .QN(n2885) );
  DFE1 \mem_reg_135][18  ( .D(D_18), .E(n6303), .C(wclk), .QN(n2886) );
  DFE1 \mem_reg_135][17  ( .D(D_17), .E(n6303), .C(wclk), .QN(n2887) );
  DFE1 \mem_reg_135][16  ( .D(D_16), .E(n6303), .C(wclk), .QN(n2888) );
  DFE1 \mem_reg_135][15  ( .D(D_15), .E(n6303), .C(wclk), .QN(n2889) );
  DFE1 \mem_reg_135][14  ( .D(D_14), .E(n6303), .C(wclk), .QN(n2890) );
  DFE1 \mem_reg_135][13  ( .D(D_13), .E(n6303), .C(wclk), .QN(n2891) );
  DFE1 \mem_reg_135][12  ( .D(D_12), .E(n6303), .C(wclk), .QN(n2892) );
  DFE1 \mem_reg_135][11  ( .D(D_11), .E(n6303), .C(wclk), .QN(n2893) );
  DFE1 \mem_reg_135][10  ( .D(D_10), .E(n6303), .C(wclk), .QN(n2894) );
  DFE1 \mem_reg_135][9  ( .D(D_9), .E(n6303), .C(wclk), .QN(n2895) );
  DFE1 \mem_reg_135][8  ( .D(D_8), .E(n6303), .C(wclk), .QN(n2896) );
  DFE1 \mem_reg_135][7  ( .D(D_7), .E(n6303), .C(wclk), .QN(n2897) );
  DFE1 \mem_reg_135][6  ( .D(D_6), .E(n6303), .C(wclk), .QN(n2898) );
  DFE1 \mem_reg_135][5  ( .D(D_5), .E(n6303), .C(wclk), .QN(n2899) );
  DFE1 \mem_reg_135][4  ( .D(D_4), .E(n6303), .C(wclk), .QN(n2900) );
  DFE1 \mem_reg_135][3  ( .D(D_3), .E(n6303), .C(wclk), .QN(n2901) );
  DFE1 \mem_reg_135][2  ( .D(D_2), .E(n6303), .C(wclk), .QN(n2902) );
  DFE1 \mem_reg_135][1  ( .D(D_1), .E(n6303), .C(wclk), .QN(n2903) );
  DFE1 \mem_reg_135][0  ( .D(D_0), .E(n6303), .C(wclk), .QN(n2904) );
  DFE1 \mem_reg_134][23  ( .D(D_23), .E(n6302), .C(wclk), .QN(n2905) );
  DFE1 \mem_reg_134][22  ( .D(D_22), .E(n6302), .C(wclk), .QN(n2906) );
  DFE1 \mem_reg_134][21  ( .D(D_21), .E(n6302), .C(wclk), .QN(n2907) );
  DFE1 \mem_reg_134][20  ( .D(D_20), .E(n6302), .C(wclk), .QN(n2908) );
  DFE1 \mem_reg_134][19  ( .D(D_19), .E(n6302), .C(wclk), .QN(n2909) );
  DFE1 \mem_reg_134][18  ( .D(D_18), .E(n6302), .C(wclk), .QN(n2910) );
  DFE1 \mem_reg_134][17  ( .D(D_17), .E(n6302), .C(wclk), .QN(n2911) );
  DFE1 \mem_reg_134][16  ( .D(D_16), .E(n6302), .C(wclk), .QN(n2912) );
  DFE1 \mem_reg_134][15  ( .D(D_15), .E(n6302), .C(wclk), .QN(n2913) );
  DFE1 \mem_reg_134][14  ( .D(D_14), .E(n6302), .C(wclk), .QN(n2914) );
  DFE1 \mem_reg_134][13  ( .D(D_13), .E(n6302), .C(wclk), .QN(n2915) );
  DFE1 \mem_reg_134][12  ( .D(D_12), .E(n6302), .C(wclk), .QN(n2916) );
  DFE1 \mem_reg_134][11  ( .D(D_11), .E(n6302), .C(wclk), .QN(n2917) );
  DFE1 \mem_reg_134][10  ( .D(D_10), .E(n6302), .C(wclk), .QN(n2918) );
  DFE1 \mem_reg_134][9  ( .D(D_9), .E(n6302), .C(wclk), .QN(n2919) );
  DFE1 \mem_reg_134][8  ( .D(D_8), .E(n6302), .C(wclk), .QN(n2920) );
  DFE1 \mem_reg_134][7  ( .D(D_7), .E(n6302), .C(wclk), .QN(n2921) );
  DFE1 \mem_reg_134][6  ( .D(D_6), .E(n6302), .C(wclk), .QN(n2922) );
  DFE1 \mem_reg_134][5  ( .D(D_5), .E(n6302), .C(wclk), .QN(n2923) );
  DFE1 \mem_reg_134][4  ( .D(D_4), .E(n6302), .C(wclk), .QN(n2924) );
  DFE1 \mem_reg_134][3  ( .D(D_3), .E(n6302), .C(wclk), .QN(n2925) );
  DFE1 \mem_reg_134][2  ( .D(D_2), .E(n6302), .C(wclk), .QN(n2926) );
  DFE1 \mem_reg_134][1  ( .D(D_1), .E(n6302), .C(wclk), .QN(n2927) );
  DFE1 \mem_reg_134][0  ( .D(D_0), .E(n6302), .C(wclk), .QN(n2928) );
  DFE1 \mem_reg_133][23  ( .D(D_23), .E(n6301), .C(wclk), .QN(n2929) );
  DFE1 \mem_reg_133][22  ( .D(D_22), .E(n6301), .C(wclk), .QN(n2930) );
  DFE1 \mem_reg_133][21  ( .D(D_21), .E(n6301), .C(wclk), .QN(n2931) );
  DFE1 \mem_reg_133][20  ( .D(D_20), .E(n6301), .C(wclk), .QN(n2932) );
  DFE1 \mem_reg_133][19  ( .D(D_19), .E(n6301), .C(wclk), .QN(n2933) );
  DFE1 \mem_reg_133][18  ( .D(D_18), .E(n6301), .C(wclk), .QN(n2934) );
  DFE1 \mem_reg_133][17  ( .D(D_17), .E(n6301), .C(wclk), .QN(n2935) );
  DFE1 \mem_reg_133][16  ( .D(D_16), .E(n6301), .C(wclk), .QN(n2936) );
  DFE1 \mem_reg_133][15  ( .D(D_15), .E(n6301), .C(wclk), .QN(n2937) );
  DFE1 \mem_reg_133][14  ( .D(D_14), .E(n6301), .C(wclk), .QN(n2938) );
  DFE1 \mem_reg_133][13  ( .D(D_13), .E(n6301), .C(wclk), .QN(n2939) );
  DFE1 \mem_reg_133][12  ( .D(D_12), .E(n6301), .C(wclk), .QN(n2940) );
  DFE1 \mem_reg_133][11  ( .D(D_11), .E(n6301), .C(wclk), .QN(n2941) );
  DFE1 \mem_reg_133][10  ( .D(D_10), .E(n6301), .C(wclk), .QN(n2942) );
  DFE1 \mem_reg_133][9  ( .D(D_9), .E(n6301), .C(wclk), .QN(n2943) );
  DFE1 \mem_reg_133][8  ( .D(D_8), .E(n6301), .C(wclk), .QN(n2944) );
  DFE1 \mem_reg_133][7  ( .D(D_7), .E(n6301), .C(wclk), .QN(n2945) );
  DFE1 \mem_reg_133][6  ( .D(D_6), .E(n6301), .C(wclk), .QN(n2946) );
  DFE1 \mem_reg_133][5  ( .D(D_5), .E(n6301), .C(wclk), .QN(n2947) );
  DFE1 \mem_reg_133][4  ( .D(D_4), .E(n6301), .C(wclk), .QN(n2948) );
  DFE1 \mem_reg_133][3  ( .D(D_3), .E(n6301), .C(wclk), .QN(n2949) );
  DFE1 \mem_reg_133][2  ( .D(D_2), .E(n6301), .C(wclk), .QN(n2950) );
  DFE1 \mem_reg_133][1  ( .D(D_1), .E(n6301), .C(wclk), .QN(n2951) );
  DFE1 \mem_reg_133][0  ( .D(D_0), .E(n6301), .C(wclk), .QN(n2952) );
  DFE1 \mem_reg_132][23  ( .D(D_23), .E(n6300), .C(wclk), .QN(n2953) );
  DFE1 \mem_reg_132][22  ( .D(D_22), .E(n6300), .C(wclk), .QN(n2954) );
  DFE1 \mem_reg_132][21  ( .D(D_21), .E(n6300), .C(wclk), .QN(n2955) );
  DFE1 \mem_reg_132][20  ( .D(D_20), .E(n6300), .C(wclk), .QN(n2956) );
  DFE1 \mem_reg_132][19  ( .D(D_19), .E(n6300), .C(wclk), .QN(n2957) );
  DFE1 \mem_reg_132][18  ( .D(D_18), .E(n6300), .C(wclk), .QN(n2958) );
  DFE1 \mem_reg_132][17  ( .D(D_17), .E(n6300), .C(wclk), .QN(n2959) );
  DFE1 \mem_reg_132][16  ( .D(D_16), .E(n6300), .C(wclk), .QN(n2960) );
  DFE1 \mem_reg_132][15  ( .D(D_15), .E(n6300), .C(wclk), .QN(n2961) );
  DFE1 \mem_reg_132][14  ( .D(D_14), .E(n6300), .C(wclk), .QN(n2962) );
  DFE1 \mem_reg_132][13  ( .D(D_13), .E(n6300), .C(wclk), .QN(n2963) );
  DFE1 \mem_reg_132][12  ( .D(D_12), .E(n6300), .C(wclk), .QN(n2964) );
  DFE1 \mem_reg_132][11  ( .D(D_11), .E(n6300), .C(wclk), .QN(n2965) );
  DFE1 \mem_reg_132][10  ( .D(D_10), .E(n6300), .C(wclk), .QN(n2966) );
  DFE1 \mem_reg_132][9  ( .D(D_9), .E(n6300), .C(wclk), .QN(n2967) );
  DFE1 \mem_reg_132][8  ( .D(D_8), .E(n6300), .C(wclk), .QN(n2968) );
  DFE1 \mem_reg_132][7  ( .D(D_7), .E(n6300), .C(wclk), .QN(n2969) );
  DFE1 \mem_reg_132][6  ( .D(D_6), .E(n6300), .C(wclk), .QN(n2970) );
  DFE1 \mem_reg_132][5  ( .D(D_5), .E(n6300), .C(wclk), .QN(n2971) );
  DFE1 \mem_reg_132][4  ( .D(D_4), .E(n6300), .C(wclk), .QN(n2972) );
  DFE1 \mem_reg_132][3  ( .D(D_3), .E(n6300), .C(wclk), .QN(n2973) );
  DFE1 \mem_reg_132][2  ( .D(D_2), .E(n6300), .C(wclk), .QN(n2974) );
  DFE1 \mem_reg_132][1  ( .D(D_1), .E(n6300), .C(wclk), .QN(n2975) );
  DFE1 \mem_reg_132][0  ( .D(D_0), .E(n6300), .C(wclk), .QN(n2976) );
  DFE1 \mem_reg_131][23  ( .D(D_23), .E(n6299), .C(wclk), .QN(n2977) );
  DFE1 \mem_reg_131][22  ( .D(D_22), .E(n6299), .C(wclk), .QN(n2978) );
  DFE1 \mem_reg_131][21  ( .D(D_21), .E(n6299), .C(wclk), .QN(n2979) );
  DFE1 \mem_reg_131][20  ( .D(D_20), .E(n6299), .C(wclk), .QN(n2980) );
  DFE1 \mem_reg_131][19  ( .D(D_19), .E(n6299), .C(wclk), .QN(n2981) );
  DFE1 \mem_reg_131][18  ( .D(D_18), .E(n6299), .C(wclk), .QN(n2982) );
  DFE1 \mem_reg_131][17  ( .D(D_17), .E(n6299), .C(wclk), .QN(n2983) );
  DFE1 \mem_reg_131][16  ( .D(D_16), .E(n6299), .C(wclk), .QN(n2984) );
  DFE1 \mem_reg_131][15  ( .D(D_15), .E(n6299), .C(wclk), .QN(n2985) );
  DFE1 \mem_reg_131][14  ( .D(D_14), .E(n6299), .C(wclk), .QN(n2986) );
  DFE1 \mem_reg_131][13  ( .D(D_13), .E(n6299), .C(wclk), .QN(n2987) );
  DFE1 \mem_reg_131][12  ( .D(D_12), .E(n6299), .C(wclk), .QN(n2988) );
  DFE1 \mem_reg_131][11  ( .D(D_11), .E(n6299), .C(wclk), .QN(n2989) );
  DFE1 \mem_reg_131][10  ( .D(D_10), .E(n6299), .C(wclk), .QN(n2990) );
  DFE1 \mem_reg_131][9  ( .D(D_9), .E(n6299), .C(wclk), .QN(n2991) );
  DFE1 \mem_reg_131][8  ( .D(D_8), .E(n6299), .C(wclk), .QN(n2992) );
  DFE1 \mem_reg_131][7  ( .D(D_7), .E(n6299), .C(wclk), .QN(n2993) );
  DFE1 \mem_reg_131][6  ( .D(D_6), .E(n6299), .C(wclk), .QN(n2994) );
  DFE1 \mem_reg_131][5  ( .D(D_5), .E(n6299), .C(wclk), .QN(n2995) );
  DFE1 \mem_reg_131][4  ( .D(D_4), .E(n6299), .C(wclk), .QN(n2996) );
  DFE1 \mem_reg_131][3  ( .D(D_3), .E(n6299), .C(wclk), .QN(n2997) );
  DFE1 \mem_reg_131][2  ( .D(D_2), .E(n6299), .C(wclk), .QN(n2998) );
  DFE1 \mem_reg_131][1  ( .D(D_1), .E(n6299), .C(wclk), .QN(n2999) );
  DFE1 \mem_reg_131][0  ( .D(D_0), .E(n6299), .C(wclk), .QN(n3000) );
  DFE1 \mem_reg_130][23  ( .D(D_23), .E(n6298), .C(wclk), .QN(n3001) );
  DFE1 \mem_reg_130][22  ( .D(D_22), .E(n6298), .C(wclk), .QN(n3002) );
  DFE1 \mem_reg_130][21  ( .D(D_21), .E(n6298), .C(wclk), .QN(n3003) );
  DFE1 \mem_reg_130][20  ( .D(D_20), .E(n6298), .C(wclk), .QN(n3004) );
  DFE1 \mem_reg_130][19  ( .D(D_19), .E(n6298), .C(wclk), .QN(n3005) );
  DFE1 \mem_reg_130][18  ( .D(D_18), .E(n6298), .C(wclk), .QN(n3006) );
  DFE1 \mem_reg_130][17  ( .D(D_17), .E(n6298), .C(wclk), .QN(n3007) );
  DFE1 \mem_reg_130][16  ( .D(D_16), .E(n6298), .C(wclk), .QN(n3008) );
  DFE1 \mem_reg_130][15  ( .D(D_15), .E(n6298), .C(wclk), .QN(n3009) );
  DFE1 \mem_reg_130][14  ( .D(D_14), .E(n6298), .C(wclk), .QN(n3010) );
  DFE1 \mem_reg_130][13  ( .D(D_13), .E(n6298), .C(wclk), .QN(n3011) );
  DFE1 \mem_reg_130][12  ( .D(D_12), .E(n6298), .C(wclk), .QN(n3012) );
  DFE1 \mem_reg_130][11  ( .D(D_11), .E(n6298), .C(wclk), .QN(n3013) );
  DFE1 \mem_reg_130][10  ( .D(D_10), .E(n6298), .C(wclk), .QN(n3014) );
  DFE1 \mem_reg_130][9  ( .D(D_9), .E(n6298), .C(wclk), .QN(n3015) );
  DFE1 \mem_reg_130][8  ( .D(D_8), .E(n6298), .C(wclk), .QN(n3016) );
  DFE1 \mem_reg_130][7  ( .D(D_7), .E(n6298), .C(wclk), .QN(n3017) );
  DFE1 \mem_reg_130][6  ( .D(D_6), .E(n6298), .C(wclk), .QN(n3018) );
  DFE1 \mem_reg_130][5  ( .D(D_5), .E(n6298), .C(wclk), .QN(n3019) );
  DFE1 \mem_reg_130][4  ( .D(D_4), .E(n6298), .C(wclk), .QN(n3020) );
  DFE1 \mem_reg_130][3  ( .D(D_3), .E(n6298), .C(wclk), .QN(n3021) );
  DFE1 \mem_reg_130][2  ( .D(D_2), .E(n6298), .C(wclk), .QN(n3022) );
  DFE1 \mem_reg_130][1  ( .D(D_1), .E(n6298), .C(wclk), .QN(n3023) );
  DFE1 \mem_reg_130][0  ( .D(D_0), .E(n6298), .C(wclk), .QN(n3024) );
  DFE1 \mem_reg_129][23  ( .D(D_23), .E(n6297), .C(wclk), .QN(n3025) );
  DFE1 \mem_reg_129][22  ( .D(D_22), .E(n6297), .C(wclk), .QN(n3026) );
  DFE1 \mem_reg_129][21  ( .D(D_21), .E(n6297), .C(wclk), .QN(n3027) );
  DFE1 \mem_reg_129][20  ( .D(D_20), .E(n6297), .C(wclk), .QN(n3028) );
  DFE1 \mem_reg_129][19  ( .D(D_19), .E(n6297), .C(wclk), .QN(n3029) );
  DFE1 \mem_reg_129][18  ( .D(D_18), .E(n6297), .C(wclk), .QN(n3030) );
  DFE1 \mem_reg_129][17  ( .D(D_17), .E(n6297), .C(wclk), .QN(n3031) );
  DFE1 \mem_reg_129][16  ( .D(D_16), .E(n6297), .C(wclk), .QN(n3032) );
  DFE1 \mem_reg_129][15  ( .D(D_15), .E(n6297), .C(wclk), .QN(n3033) );
  DFE1 \mem_reg_129][14  ( .D(D_14), .E(n6297), .C(wclk), .QN(n3034) );
  DFE1 \mem_reg_129][13  ( .D(D_13), .E(n6297), .C(wclk), .QN(n3035) );
  DFE1 \mem_reg_129][12  ( .D(D_12), .E(n6297), .C(wclk), .QN(n3036) );
  DFE1 \mem_reg_129][11  ( .D(D_11), .E(n6297), .C(wclk), .QN(n3037) );
  DFE1 \mem_reg_129][10  ( .D(D_10), .E(n6297), .C(wclk), .QN(n3038) );
  DFE1 \mem_reg_129][9  ( .D(D_9), .E(n6297), .C(wclk), .QN(n3039) );
  DFE1 \mem_reg_129][8  ( .D(D_8), .E(n6297), .C(wclk), .QN(n3040) );
  DFE1 \mem_reg_129][7  ( .D(D_7), .E(n6297), .C(wclk), .QN(n3041) );
  DFE1 \mem_reg_129][6  ( .D(D_6), .E(n6297), .C(wclk), .QN(n3042) );
  DFE1 \mem_reg_129][5  ( .D(D_5), .E(n6297), .C(wclk), .QN(n3043) );
  DFE1 \mem_reg_129][4  ( .D(D_4), .E(n6297), .C(wclk), .QN(n3044) );
  DFE1 \mem_reg_129][3  ( .D(D_3), .E(n6297), .C(wclk), .QN(n3045) );
  DFE1 \mem_reg_129][2  ( .D(D_2), .E(n6297), .C(wclk), .QN(n3046) );
  DFE1 \mem_reg_129][1  ( .D(D_1), .E(n6297), .C(wclk), .QN(n3047) );
  DFE1 \mem_reg_129][0  ( .D(D_0), .E(n6297), .C(wclk), .QN(n3048) );
  DFE1 \mem_reg_128][23  ( .D(D_23), .E(n6295), .C(wclk), .QN(n3049) );
  DFE1 \mem_reg_128][22  ( .D(D_22), .E(n6295), .C(wclk), .QN(n3050) );
  DFE1 \mem_reg_128][21  ( .D(D_21), .E(n6295), .C(wclk), .QN(n3051) );
  DFE1 \mem_reg_128][20  ( .D(D_20), .E(n6295), .C(wclk), .QN(n3052) );
  DFE1 \mem_reg_128][19  ( .D(D_19), .E(n6295), .C(wclk), .QN(n3053) );
  DFE1 \mem_reg_128][18  ( .D(D_18), .E(n6295), .C(wclk), .QN(n3054) );
  DFE1 \mem_reg_128][17  ( .D(D_17), .E(n6295), .C(wclk), .QN(n3055) );
  DFE1 \mem_reg_128][16  ( .D(D_16), .E(n6295), .C(wclk), .QN(n3056) );
  DFE1 \mem_reg_128][15  ( .D(D_15), .E(n6295), .C(wclk), .QN(n3057) );
  DFE1 \mem_reg_128][14  ( .D(D_14), .E(n6295), .C(wclk), .QN(n3058) );
  DFE1 \mem_reg_128][13  ( .D(D_13), .E(n6295), .C(wclk), .QN(n3059) );
  DFE1 \mem_reg_128][12  ( .D(D_12), .E(n6295), .C(wclk), .QN(n3060) );
  DFE1 \mem_reg_128][11  ( .D(D_11), .E(n6295), .C(wclk), .QN(n3061) );
  DFE1 \mem_reg_128][10  ( .D(D_10), .E(n6295), .C(wclk), .QN(n3062) );
  DFE1 \mem_reg_128][9  ( .D(D_9), .E(n6295), .C(wclk), .QN(n3063) );
  DFE1 \mem_reg_128][8  ( .D(D_8), .E(n6295), .C(wclk), .QN(n3064) );
  DFE1 \mem_reg_128][7  ( .D(D_7), .E(n6295), .C(wclk), .QN(n3065) );
  DFE1 \mem_reg_128][6  ( .D(D_6), .E(n6295), .C(wclk), .QN(n3066) );
  DFE1 \mem_reg_128][5  ( .D(D_5), .E(n6295), .C(wclk), .QN(n3067) );
  DFE1 \mem_reg_128][4  ( .D(D_4), .E(n6295), .C(wclk), .QN(n3068) );
  DFE1 \mem_reg_128][3  ( .D(D_3), .E(n6295), .C(wclk), .QN(n3069) );
  DFE1 \mem_reg_128][2  ( .D(D_2), .E(n6295), .C(wclk), .QN(n3070) );
  DFE1 \mem_reg_128][1  ( .D(D_1), .E(n6295), .C(wclk), .QN(n3071) );
  DFE1 \mem_reg_128][0  ( .D(D_0), .E(n6295), .C(wclk), .QN(n3072) );
  DFE1 \mem_reg_127][23  ( .D(D_23), .E(n6293), .C(wclk), .QN(n3073) );
  DFE1 \mem_reg_127][22  ( .D(D_22), .E(n6293), .C(wclk), .QN(n3074) );
  DFE1 \mem_reg_127][21  ( .D(D_21), .E(n6293), .C(wclk), .QN(n3075) );
  DFE1 \mem_reg_127][20  ( .D(D_20), .E(n6293), .C(wclk), .QN(n3076) );
  DFE1 \mem_reg_127][19  ( .D(D_19), .E(n6293), .C(wclk), .QN(n3077) );
  DFE1 \mem_reg_127][18  ( .D(D_18), .E(n6293), .C(wclk), .QN(n3078) );
  DFE1 \mem_reg_127][17  ( .D(D_17), .E(n6293), .C(wclk), .QN(n3079) );
  DFE1 \mem_reg_127][16  ( .D(D_16), .E(n6293), .C(wclk), .QN(n3080) );
  DFE1 \mem_reg_127][15  ( .D(D_15), .E(n6293), .C(wclk), .QN(n3081) );
  DFE1 \mem_reg_127][14  ( .D(D_14), .E(n6293), .C(wclk), .QN(n3082) );
  DFE1 \mem_reg_127][13  ( .D(D_13), .E(n6293), .C(wclk), .QN(n3083) );
  DFE1 \mem_reg_127][12  ( .D(D_12), .E(n6293), .C(wclk), .QN(n3084) );
  DFE1 \mem_reg_127][11  ( .D(D_11), .E(n6293), .C(wclk), .QN(n3085) );
  DFE1 \mem_reg_127][10  ( .D(D_10), .E(n6293), .C(wclk), .QN(n3086) );
  DFE1 \mem_reg_127][9  ( .D(D_9), .E(n6293), .C(wclk), .QN(n3087) );
  DFE1 \mem_reg_127][8  ( .D(D_8), .E(n6293), .C(wclk), .QN(n3088) );
  DFE1 \mem_reg_127][7  ( .D(D_7), .E(n6293), .C(wclk), .QN(n3089) );
  DFE1 \mem_reg_127][6  ( .D(D_6), .E(n6293), .C(wclk), .QN(n3090) );
  DFE1 \mem_reg_127][5  ( .D(D_5), .E(n6293), .C(wclk), .QN(n3091) );
  DFE1 \mem_reg_127][4  ( .D(D_4), .E(n6293), .C(wclk), .QN(n3092) );
  DFE1 \mem_reg_127][3  ( .D(D_3), .E(n6293), .C(wclk), .QN(n3093) );
  DFE1 \mem_reg_127][2  ( .D(D_2), .E(n6293), .C(wclk), .QN(n3094) );
  DFE1 \mem_reg_127][1  ( .D(D_1), .E(n6293), .C(wclk), .QN(n3095) );
  DFE1 \mem_reg_127][0  ( .D(D_0), .E(n6293), .C(wclk), .QN(n3096) );
  DFE1 \mem_reg_126][23  ( .D(D_23), .E(n6292), .C(wclk), .QN(n3097) );
  DFE1 \mem_reg_126][22  ( .D(D_22), .E(n6292), .C(wclk), .QN(n3098) );
  DFE1 \mem_reg_126][21  ( .D(D_21), .E(n6292), .C(wclk), .QN(n3099) );
  DFE1 \mem_reg_126][20  ( .D(D_20), .E(n6292), .C(wclk), .QN(n3100) );
  DFE1 \mem_reg_126][19  ( .D(D_19), .E(n6292), .C(wclk), .QN(n3101) );
  DFE1 \mem_reg_126][18  ( .D(D_18), .E(n6292), .C(wclk), .QN(n3102) );
  DFE1 \mem_reg_126][17  ( .D(D_17), .E(n6292), .C(wclk), .QN(n3103) );
  DFE1 \mem_reg_126][16  ( .D(D_16), .E(n6292), .C(wclk), .QN(n3104) );
  DFE1 \mem_reg_126][15  ( .D(D_15), .E(n6292), .C(wclk), .QN(n3105) );
  DFE1 \mem_reg_126][14  ( .D(D_14), .E(n6292), .C(wclk), .QN(n3106) );
  DFE1 \mem_reg_126][13  ( .D(D_13), .E(n6292), .C(wclk), .QN(n3107) );
  DFE1 \mem_reg_126][12  ( .D(D_12), .E(n6292), .C(wclk), .QN(n3108) );
  DFE1 \mem_reg_126][11  ( .D(D_11), .E(n6292), .C(wclk), .QN(n3109) );
  DFE1 \mem_reg_126][10  ( .D(D_10), .E(n6292), .C(wclk), .QN(n3110) );
  DFE1 \mem_reg_126][9  ( .D(D_9), .E(n6292), .C(wclk), .QN(n3111) );
  DFE1 \mem_reg_126][8  ( .D(D_8), .E(n6292), .C(wclk), .QN(n3112) );
  DFE1 \mem_reg_126][7  ( .D(D_7), .E(n6292), .C(wclk), .QN(n3113) );
  DFE1 \mem_reg_126][6  ( .D(D_6), .E(n6292), .C(wclk), .QN(n3114) );
  DFE1 \mem_reg_126][5  ( .D(D_5), .E(n6292), .C(wclk), .QN(n3115) );
  DFE1 \mem_reg_126][4  ( .D(D_4), .E(n6292), .C(wclk), .QN(n3116) );
  DFE1 \mem_reg_126][3  ( .D(D_3), .E(n6292), .C(wclk), .QN(n3117) );
  DFE1 \mem_reg_126][2  ( .D(D_2), .E(n6292), .C(wclk), .QN(n3118) );
  DFE1 \mem_reg_126][1  ( .D(D_1), .E(n6292), .C(wclk), .QN(n3119) );
  DFE1 \mem_reg_126][0  ( .D(D_0), .E(n6292), .C(wclk), .QN(n3120) );
  DFE1 \mem_reg_125][23  ( .D(D_23), .E(n6291), .C(wclk), .QN(n3121) );
  DFE1 \mem_reg_125][22  ( .D(D_22), .E(n6291), .C(wclk), .QN(n3122) );
  DFE1 \mem_reg_125][21  ( .D(D_21), .E(n6291), .C(wclk), .QN(n3123) );
  DFE1 \mem_reg_125][20  ( .D(D_20), .E(n6291), .C(wclk), .QN(n3124) );
  DFE1 \mem_reg_125][19  ( .D(D_19), .E(n6291), .C(wclk), .QN(n3125) );
  DFE1 \mem_reg_125][18  ( .D(D_18), .E(n6291), .C(wclk), .QN(n3126) );
  DFE1 \mem_reg_125][17  ( .D(D_17), .E(n6291), .C(wclk), .QN(n3127) );
  DFE1 \mem_reg_125][16  ( .D(D_16), .E(n6291), .C(wclk), .QN(n3128) );
  DFE1 \mem_reg_125][15  ( .D(D_15), .E(n6291), .C(wclk), .QN(n3129) );
  DFE1 \mem_reg_125][14  ( .D(D_14), .E(n6291), .C(wclk), .QN(n3130) );
  DFE1 \mem_reg_125][13  ( .D(D_13), .E(n6291), .C(wclk), .QN(n3131) );
  DFE1 \mem_reg_125][12  ( .D(D_12), .E(n6291), .C(wclk), .QN(n3132) );
  DFE1 \mem_reg_125][11  ( .D(D_11), .E(n6291), .C(wclk), .QN(n3133) );
  DFE1 \mem_reg_125][10  ( .D(D_10), .E(n6291), .C(wclk), .QN(n3134) );
  DFE1 \mem_reg_125][9  ( .D(D_9), .E(n6291), .C(wclk), .QN(n3135) );
  DFE1 \mem_reg_125][8  ( .D(D_8), .E(n6291), .C(wclk), .QN(n3136) );
  DFE1 \mem_reg_125][7  ( .D(D_7), .E(n6291), .C(wclk), .QN(n3137) );
  DFE1 \mem_reg_125][6  ( .D(D_6), .E(n6291), .C(wclk), .QN(n3138) );
  DFE1 \mem_reg_125][5  ( .D(D_5), .E(n6291), .C(wclk), .QN(n3139) );
  DFE1 \mem_reg_125][4  ( .D(D_4), .E(n6291), .C(wclk), .QN(n3140) );
  DFE1 \mem_reg_125][3  ( .D(D_3), .E(n6291), .C(wclk), .QN(n3141) );
  DFE1 \mem_reg_125][2  ( .D(D_2), .E(n6291), .C(wclk), .QN(n3142) );
  DFE1 \mem_reg_125][1  ( .D(D_1), .E(n6291), .C(wclk), .QN(n3143) );
  DFE1 \mem_reg_125][0  ( .D(D_0), .E(n6291), .C(wclk), .QN(n3144) );
  DFE1 \mem_reg_124][23  ( .D(D_23), .E(n6290), .C(wclk), .QN(n3145) );
  DFE1 \mem_reg_124][22  ( .D(D_22), .E(n6290), .C(wclk), .QN(n3146) );
  DFE1 \mem_reg_124][21  ( .D(D_21), .E(n6290), .C(wclk), .QN(n3147) );
  DFE1 \mem_reg_124][20  ( .D(D_20), .E(n6290), .C(wclk), .QN(n3148) );
  DFE1 \mem_reg_124][19  ( .D(D_19), .E(n6290), .C(wclk), .QN(n3149) );
  DFE1 \mem_reg_124][18  ( .D(D_18), .E(n6290), .C(wclk), .QN(n3150) );
  DFE1 \mem_reg_124][17  ( .D(D_17), .E(n6290), .C(wclk), .QN(n3151) );
  DFE1 \mem_reg_124][16  ( .D(D_16), .E(n6290), .C(wclk), .QN(n3152) );
  DFE1 \mem_reg_124][15  ( .D(D_15), .E(n6290), .C(wclk), .QN(n3153) );
  DFE1 \mem_reg_124][14  ( .D(D_14), .E(n6290), .C(wclk), .QN(n3154) );
  DFE1 \mem_reg_124][13  ( .D(D_13), .E(n6290), .C(wclk), .QN(n3155) );
  DFE1 \mem_reg_124][12  ( .D(D_12), .E(n6290), .C(wclk), .QN(n3156) );
  DFE1 \mem_reg_124][11  ( .D(D_11), .E(n6290), .C(wclk), .QN(n3157) );
  DFE1 \mem_reg_124][10  ( .D(D_10), .E(n6290), .C(wclk), .QN(n3158) );
  DFE1 \mem_reg_124][9  ( .D(D_9), .E(n6290), .C(wclk), .QN(n3159) );
  DFE1 \mem_reg_124][8  ( .D(D_8), .E(n6290), .C(wclk), .QN(n3160) );
  DFE1 \mem_reg_124][7  ( .D(D_7), .E(n6290), .C(wclk), .QN(n3161) );
  DFE1 \mem_reg_124][6  ( .D(D_6), .E(n6290), .C(wclk), .QN(n3162) );
  DFE1 \mem_reg_124][5  ( .D(D_5), .E(n6290), .C(wclk), .QN(n3163) );
  DFE1 \mem_reg_124][4  ( .D(D_4), .E(n6290), .C(wclk), .QN(n3164) );
  DFE1 \mem_reg_124][3  ( .D(D_3), .E(n6290), .C(wclk), .QN(n3165) );
  DFE1 \mem_reg_124][2  ( .D(D_2), .E(n6290), .C(wclk), .QN(n3166) );
  DFE1 \mem_reg_124][1  ( .D(D_1), .E(n6290), .C(wclk), .QN(n3167) );
  DFE1 \mem_reg_124][0  ( .D(D_0), .E(n6290), .C(wclk), .QN(n3168) );
  DFE1 \mem_reg_123][23  ( .D(D_23), .E(n6288), .C(wclk), .QN(n3169) );
  DFE1 \mem_reg_123][22  ( .D(D_22), .E(n6288), .C(wclk), .QN(n3170) );
  DFE1 \mem_reg_123][21  ( .D(D_21), .E(n6288), .C(wclk), .QN(n3171) );
  DFE1 \mem_reg_123][20  ( .D(D_20), .E(n6288), .C(wclk), .QN(n3172) );
  DFE1 \mem_reg_123][19  ( .D(D_19), .E(n6288), .C(wclk), .QN(n3173) );
  DFE1 \mem_reg_123][18  ( .D(D_18), .E(n6288), .C(wclk), .QN(n3174) );
  DFE1 \mem_reg_123][17  ( .D(D_17), .E(n6288), .C(wclk), .QN(n3175) );
  DFE1 \mem_reg_123][16  ( .D(D_16), .E(n6288), .C(wclk), .QN(n3176) );
  DFE1 \mem_reg_123][15  ( .D(D_15), .E(n6288), .C(wclk), .QN(n3177) );
  DFE1 \mem_reg_123][14  ( .D(D_14), .E(n6288), .C(wclk), .QN(n3178) );
  DFE1 \mem_reg_123][13  ( .D(D_13), .E(n6288), .C(wclk), .QN(n3179) );
  DFE1 \mem_reg_123][12  ( .D(D_12), .E(n6288), .C(wclk), .QN(n3180) );
  DFE1 \mem_reg_123][11  ( .D(D_11), .E(n6288), .C(wclk), .QN(n3181) );
  DFE1 \mem_reg_123][10  ( .D(D_10), .E(n6288), .C(wclk), .QN(n3182) );
  DFE1 \mem_reg_123][9  ( .D(D_9), .E(n6288), .C(wclk), .QN(n3183) );
  DFE1 \mem_reg_123][8  ( .D(D_8), .E(n6288), .C(wclk), .QN(n3184) );
  DFE1 \mem_reg_123][7  ( .D(D_7), .E(n6288), .C(wclk), .QN(n3185) );
  DFE1 \mem_reg_123][6  ( .D(D_6), .E(n6288), .C(wclk), .QN(n3186) );
  DFE1 \mem_reg_123][5  ( .D(D_5), .E(n6288), .C(wclk), .QN(n3187) );
  DFE1 \mem_reg_123][4  ( .D(D_4), .E(n6288), .C(wclk), .QN(n3188) );
  DFE1 \mem_reg_123][3  ( .D(D_3), .E(n6288), .C(wclk), .QN(n3189) );
  DFE1 \mem_reg_123][2  ( .D(D_2), .E(n6288), .C(wclk), .QN(n3190) );
  DFE1 \mem_reg_123][1  ( .D(D_1), .E(n6288), .C(wclk), .QN(n3191) );
  DFE1 \mem_reg_123][0  ( .D(D_0), .E(n6288), .C(wclk), .QN(n3192) );
  DFE1 \mem_reg_122][23  ( .D(D_23), .E(n6287), .C(wclk), .QN(n3193) );
  DFE1 \mem_reg_122][22  ( .D(D_22), .E(n6287), .C(wclk), .QN(n3194) );
  DFE1 \mem_reg_122][21  ( .D(D_21), .E(n6287), .C(wclk), .QN(n3195) );
  DFE1 \mem_reg_122][20  ( .D(D_20), .E(n6287), .C(wclk), .QN(n3196) );
  DFE1 \mem_reg_122][19  ( .D(D_19), .E(n6287), .C(wclk), .QN(n3197) );
  DFE1 \mem_reg_122][18  ( .D(D_18), .E(n6287), .C(wclk), .QN(n3198) );
  DFE1 \mem_reg_122][17  ( .D(D_17), .E(n6287), .C(wclk), .QN(n3199) );
  DFE1 \mem_reg_122][16  ( .D(D_16), .E(n6287), .C(wclk), .QN(n3200) );
  DFE1 \mem_reg_122][15  ( .D(D_15), .E(n6287), .C(wclk), .QN(n3201) );
  DFE1 \mem_reg_122][14  ( .D(D_14), .E(n6287), .C(wclk), .QN(n3202) );
  DFE1 \mem_reg_122][13  ( .D(D_13), .E(n6287), .C(wclk), .QN(n3203) );
  DFE1 \mem_reg_122][12  ( .D(D_12), .E(n6287), .C(wclk), .QN(n3204) );
  DFE1 \mem_reg_122][11  ( .D(D_11), .E(n6287), .C(wclk), .QN(n3205) );
  DFE1 \mem_reg_122][10  ( .D(D_10), .E(n6287), .C(wclk), .QN(n3206) );
  DFE1 \mem_reg_122][9  ( .D(D_9), .E(n6287), .C(wclk), .QN(n3207) );
  DFE1 \mem_reg_122][8  ( .D(D_8), .E(n6287), .C(wclk), .QN(n3208) );
  DFE1 \mem_reg_122][7  ( .D(D_7), .E(n6287), .C(wclk), .QN(n3209) );
  DFE1 \mem_reg_122][6  ( .D(D_6), .E(n6287), .C(wclk), .QN(n3210) );
  DFE1 \mem_reg_122][5  ( .D(D_5), .E(n6287), .C(wclk), .QN(n3211) );
  DFE1 \mem_reg_122][4  ( .D(D_4), .E(n6287), .C(wclk), .QN(n3212) );
  DFE1 \mem_reg_122][3  ( .D(D_3), .E(n6287), .C(wclk), .QN(n3213) );
  DFE1 \mem_reg_122][2  ( .D(D_2), .E(n6287), .C(wclk), .QN(n3214) );
  DFE1 \mem_reg_122][1  ( .D(D_1), .E(n6287), .C(wclk), .QN(n3215) );
  DFE1 \mem_reg_122][0  ( .D(D_0), .E(n6287), .C(wclk), .QN(n3216) );
  DFE1 \mem_reg_121][23  ( .D(D_23), .E(n6286), .C(wclk), .QN(n3217) );
  DFE1 \mem_reg_121][22  ( .D(D_22), .E(n6286), .C(wclk), .QN(n3218) );
  DFE1 \mem_reg_121][21  ( .D(D_21), .E(n6286), .C(wclk), .QN(n3219) );
  DFE1 \mem_reg_121][20  ( .D(D_20), .E(n6286), .C(wclk), .QN(n3220) );
  DFE1 \mem_reg_121][19  ( .D(D_19), .E(n6286), .C(wclk), .QN(n3221) );
  DFE1 \mem_reg_121][18  ( .D(D_18), .E(n6286), .C(wclk), .QN(n3222) );
  DFE1 \mem_reg_121][17  ( .D(D_17), .E(n6286), .C(wclk), .QN(n3223) );
  DFE1 \mem_reg_121][16  ( .D(D_16), .E(n6286), .C(wclk), .QN(n3224) );
  DFE1 \mem_reg_121][15  ( .D(D_15), .E(n6286), .C(wclk), .QN(n3225) );
  DFE1 \mem_reg_121][14  ( .D(D_14), .E(n6286), .C(wclk), .QN(n3226) );
  DFE1 \mem_reg_121][13  ( .D(D_13), .E(n6286), .C(wclk), .QN(n3227) );
  DFE1 \mem_reg_121][12  ( .D(D_12), .E(n6286), .C(wclk), .QN(n3228) );
  DFE1 \mem_reg_121][11  ( .D(D_11), .E(n6286), .C(wclk), .QN(n3229) );
  DFE1 \mem_reg_121][10  ( .D(D_10), .E(n6286), .C(wclk), .QN(n3230) );
  DFE1 \mem_reg_121][9  ( .D(D_9), .E(n6286), .C(wclk), .QN(n3231) );
  DFE1 \mem_reg_121][8  ( .D(D_8), .E(n6286), .C(wclk), .QN(n3232) );
  DFE1 \mem_reg_121][7  ( .D(D_7), .E(n6286), .C(wclk), .QN(n3233) );
  DFE1 \mem_reg_121][6  ( .D(D_6), .E(n6286), .C(wclk), .QN(n3234) );
  DFE1 \mem_reg_121][5  ( .D(D_5), .E(n6286), .C(wclk), .QN(n3235) );
  DFE1 \mem_reg_121][4  ( .D(D_4), .E(n6286), .C(wclk), .QN(n3236) );
  DFE1 \mem_reg_121][3  ( .D(D_3), .E(n6286), .C(wclk), .QN(n3237) );
  DFE1 \mem_reg_121][2  ( .D(D_2), .E(n6286), .C(wclk), .QN(n3238) );
  DFE1 \mem_reg_121][1  ( .D(D_1), .E(n6286), .C(wclk), .QN(n3239) );
  DFE1 \mem_reg_121][0  ( .D(D_0), .E(n6286), .C(wclk), .QN(n3240) );
  DFE1 \mem_reg_120][23  ( .D(D_23), .E(n6285), .C(wclk), .QN(n3241) );
  DFE1 \mem_reg_120][22  ( .D(D_22), .E(n6285), .C(wclk), .QN(n3242) );
  DFE1 \mem_reg_120][21  ( .D(D_21), .E(n6285), .C(wclk), .QN(n3243) );
  DFE1 \mem_reg_120][20  ( .D(D_20), .E(n6285), .C(wclk), .QN(n3244) );
  DFE1 \mem_reg_120][19  ( .D(D_19), .E(n6285), .C(wclk), .QN(n3245) );
  DFE1 \mem_reg_120][18  ( .D(D_18), .E(n6285), .C(wclk), .QN(n3246) );
  DFE1 \mem_reg_120][17  ( .D(D_17), .E(n6285), .C(wclk), .QN(n3247) );
  DFE1 \mem_reg_120][16  ( .D(D_16), .E(n6285), .C(wclk), .QN(n3248) );
  DFE1 \mem_reg_120][15  ( .D(D_15), .E(n6285), .C(wclk), .QN(n3249) );
  DFE1 \mem_reg_120][14  ( .D(D_14), .E(n6285), .C(wclk), .QN(n3250) );
  DFE1 \mem_reg_120][13  ( .D(D_13), .E(n6285), .C(wclk), .QN(n3251) );
  DFE1 \mem_reg_120][12  ( .D(D_12), .E(n6285), .C(wclk), .QN(n3252) );
  DFE1 \mem_reg_120][11  ( .D(D_11), .E(n6285), .C(wclk), .QN(n3253) );
  DFE1 \mem_reg_120][10  ( .D(D_10), .E(n6285), .C(wclk), .QN(n3254) );
  DFE1 \mem_reg_120][9  ( .D(D_9), .E(n6285), .C(wclk), .QN(n3255) );
  DFE1 \mem_reg_120][8  ( .D(D_8), .E(n6285), .C(wclk), .QN(n3256) );
  DFE1 \mem_reg_120][7  ( .D(D_7), .E(n6285), .C(wclk), .QN(n3257) );
  DFE1 \mem_reg_120][6  ( .D(D_6), .E(n6285), .C(wclk), .QN(n3258) );
  DFE1 \mem_reg_120][5  ( .D(D_5), .E(n6285), .C(wclk), .QN(n3259) );
  DFE1 \mem_reg_120][4  ( .D(D_4), .E(n6285), .C(wclk), .QN(n3260) );
  DFE1 \mem_reg_120][3  ( .D(D_3), .E(n6285), .C(wclk), .QN(n3261) );
  DFE1 \mem_reg_120][2  ( .D(D_2), .E(n6285), .C(wclk), .QN(n3262) );
  DFE1 \mem_reg_120][1  ( .D(D_1), .E(n6285), .C(wclk), .QN(n3263) );
  DFE1 \mem_reg_120][0  ( .D(D_0), .E(n6285), .C(wclk), .QN(n3264) );
  DFE1 \mem_reg_119][23  ( .D(D_23), .E(n6284), .C(wclk), .QN(n3265) );
  DFE1 \mem_reg_119][22  ( .D(D_22), .E(n6284), .C(wclk), .QN(n3266) );
  DFE1 \mem_reg_119][21  ( .D(D_21), .E(n6284), .C(wclk), .QN(n3267) );
  DFE1 \mem_reg_119][20  ( .D(D_20), .E(n6284), .C(wclk), .QN(n3268) );
  DFE1 \mem_reg_119][19  ( .D(D_19), .E(n6284), .C(wclk), .QN(n3269) );
  DFE1 \mem_reg_119][18  ( .D(D_18), .E(n6284), .C(wclk), .QN(n3270) );
  DFE1 \mem_reg_119][17  ( .D(D_17), .E(n6284), .C(wclk), .QN(n3271) );
  DFE1 \mem_reg_119][16  ( .D(D_16), .E(n6284), .C(wclk), .QN(n3272) );
  DFE1 \mem_reg_119][15  ( .D(D_15), .E(n6284), .C(wclk), .QN(n3273) );
  DFE1 \mem_reg_119][14  ( .D(D_14), .E(n6284), .C(wclk), .QN(n3274) );
  DFE1 \mem_reg_119][13  ( .D(D_13), .E(n6284), .C(wclk), .QN(n3275) );
  DFE1 \mem_reg_119][12  ( .D(D_12), .E(n6284), .C(wclk), .QN(n3276) );
  DFE1 \mem_reg_119][11  ( .D(D_11), .E(n6284), .C(wclk), .QN(n3277) );
  DFE1 \mem_reg_119][10  ( .D(D_10), .E(n6284), .C(wclk), .QN(n3278) );
  DFE1 \mem_reg_119][9  ( .D(D_9), .E(n6284), .C(wclk), .QN(n3279) );
  DFE1 \mem_reg_119][8  ( .D(D_8), .E(n6284), .C(wclk), .QN(n3280) );
  DFE1 \mem_reg_119][7  ( .D(D_7), .E(n6284), .C(wclk), .QN(n3281) );
  DFE1 \mem_reg_119][6  ( .D(D_6), .E(n6284), .C(wclk), .QN(n3282) );
  DFE1 \mem_reg_119][5  ( .D(D_5), .E(n6284), .C(wclk), .QN(n3283) );
  DFE1 \mem_reg_119][4  ( .D(D_4), .E(n6284), .C(wclk), .QN(n3284) );
  DFE1 \mem_reg_119][3  ( .D(D_3), .E(n6284), .C(wclk), .QN(n3285) );
  DFE1 \mem_reg_119][2  ( .D(D_2), .E(n6284), .C(wclk), .QN(n3286) );
  DFE1 \mem_reg_119][1  ( .D(D_1), .E(n6284), .C(wclk), .QN(n3287) );
  DFE1 \mem_reg_119][0  ( .D(D_0), .E(n6284), .C(wclk), .QN(n3288) );
  DFE1 \mem_reg_118][23  ( .D(D_23), .E(n6283), .C(wclk), .QN(n3289) );
  DFE1 \mem_reg_118][22  ( .D(D_22), .E(n6283), .C(wclk), .QN(n3290) );
  DFE1 \mem_reg_118][21  ( .D(D_21), .E(n6283), .C(wclk), .QN(n3291) );
  DFE1 \mem_reg_118][20  ( .D(D_20), .E(n6283), .C(wclk), .QN(n3292) );
  DFE1 \mem_reg_118][19  ( .D(D_19), .E(n6283), .C(wclk), .QN(n3293) );
  DFE1 \mem_reg_118][18  ( .D(D_18), .E(n6283), .C(wclk), .QN(n3294) );
  DFE1 \mem_reg_118][17  ( .D(D_17), .E(n6283), .C(wclk), .QN(n3295) );
  DFE1 \mem_reg_118][16  ( .D(D_16), .E(n6283), .C(wclk), .QN(n3296) );
  DFE1 \mem_reg_118][15  ( .D(D_15), .E(n6283), .C(wclk), .QN(n3297) );
  DFE1 \mem_reg_118][14  ( .D(D_14), .E(n6283), .C(wclk), .QN(n3298) );
  DFE1 \mem_reg_118][13  ( .D(D_13), .E(n6283), .C(wclk), .QN(n3299) );
  DFE1 \mem_reg_118][12  ( .D(D_12), .E(n6283), .C(wclk), .QN(n3300) );
  DFE1 \mem_reg_118][11  ( .D(D_11), .E(n6283), .C(wclk), .QN(n3301) );
  DFE1 \mem_reg_118][10  ( .D(D_10), .E(n6283), .C(wclk), .QN(n3302) );
  DFE1 \mem_reg_118][9  ( .D(D_9), .E(n6283), .C(wclk), .QN(n3303) );
  DFE1 \mem_reg_118][8  ( .D(D_8), .E(n6283), .C(wclk), .QN(n3304) );
  DFE1 \mem_reg_118][7  ( .D(D_7), .E(n6283), .C(wclk), .QN(n3305) );
  DFE1 \mem_reg_118][6  ( .D(D_6), .E(n6283), .C(wclk), .QN(n3306) );
  DFE1 \mem_reg_118][5  ( .D(D_5), .E(n6283), .C(wclk), .QN(n3307) );
  DFE1 \mem_reg_118][4  ( .D(D_4), .E(n6283), .C(wclk), .QN(n3308) );
  DFE1 \mem_reg_118][3  ( .D(D_3), .E(n6283), .C(wclk), .QN(n3309) );
  DFE1 \mem_reg_118][2  ( .D(D_2), .E(n6283), .C(wclk), .QN(n3310) );
  DFE1 \mem_reg_118][1  ( .D(D_1), .E(n6283), .C(wclk), .QN(n3311) );
  DFE1 \mem_reg_118][0  ( .D(D_0), .E(n6283), .C(wclk), .QN(n3312) );
  DFE1 \mem_reg_117][23  ( .D(D_23), .E(n6282), .C(wclk), .QN(n3313) );
  DFE1 \mem_reg_117][22  ( .D(D_22), .E(n6282), .C(wclk), .QN(n3314) );
  DFE1 \mem_reg_117][21  ( .D(D_21), .E(n6282), .C(wclk), .QN(n3315) );
  DFE1 \mem_reg_117][20  ( .D(D_20), .E(n6282), .C(wclk), .QN(n3316) );
  DFE1 \mem_reg_117][19  ( .D(D_19), .E(n6282), .C(wclk), .QN(n3317) );
  DFE1 \mem_reg_117][18  ( .D(D_18), .E(n6282), .C(wclk), .QN(n3318) );
  DFE1 \mem_reg_117][17  ( .D(D_17), .E(n6282), .C(wclk), .QN(n3319) );
  DFE1 \mem_reg_117][16  ( .D(D_16), .E(n6282), .C(wclk), .QN(n3320) );
  DFE1 \mem_reg_117][15  ( .D(D_15), .E(n6282), .C(wclk), .QN(n3321) );
  DFE1 \mem_reg_117][14  ( .D(D_14), .E(n6282), .C(wclk), .QN(n3322) );
  DFE1 \mem_reg_117][13  ( .D(D_13), .E(n6282), .C(wclk), .QN(n3323) );
  DFE1 \mem_reg_117][12  ( .D(D_12), .E(n6282), .C(wclk), .QN(n3324) );
  DFE1 \mem_reg_117][11  ( .D(D_11), .E(n6282), .C(wclk), .QN(n3325) );
  DFE1 \mem_reg_117][10  ( .D(D_10), .E(n6282), .C(wclk), .QN(n3326) );
  DFE1 \mem_reg_117][9  ( .D(D_9), .E(n6282), .C(wclk), .QN(n3327) );
  DFE1 \mem_reg_117][8  ( .D(D_8), .E(n6282), .C(wclk), .QN(n3328) );
  DFE1 \mem_reg_117][7  ( .D(D_7), .E(n6282), .C(wclk), .QN(n3329) );
  DFE1 \mem_reg_117][6  ( .D(D_6), .E(n6282), .C(wclk), .QN(n3330) );
  DFE1 \mem_reg_117][5  ( .D(D_5), .E(n6282), .C(wclk), .QN(n3331) );
  DFE1 \mem_reg_117][4  ( .D(D_4), .E(n6282), .C(wclk), .QN(n3332) );
  DFE1 \mem_reg_117][3  ( .D(D_3), .E(n6282), .C(wclk), .QN(n3333) );
  DFE1 \mem_reg_117][2  ( .D(D_2), .E(n6282), .C(wclk), .QN(n3334) );
  DFE1 \mem_reg_117][1  ( .D(D_1), .E(n6282), .C(wclk), .QN(n3335) );
  DFE1 \mem_reg_117][0  ( .D(D_0), .E(n6282), .C(wclk), .QN(n3336) );
  DFE1 \mem_reg_116][23  ( .D(D_23), .E(n6281), .C(wclk), .QN(n3337) );
  DFE1 \mem_reg_116][22  ( .D(D_22), .E(n6281), .C(wclk), .QN(n3338) );
  DFE1 \mem_reg_116][21  ( .D(D_21), .E(n6281), .C(wclk), .QN(n3339) );
  DFE1 \mem_reg_116][20  ( .D(D_20), .E(n6281), .C(wclk), .QN(n3340) );
  DFE1 \mem_reg_116][19  ( .D(D_19), .E(n6281), .C(wclk), .QN(n3341) );
  DFE1 \mem_reg_116][18  ( .D(D_18), .E(n6281), .C(wclk), .QN(n3342) );
  DFE1 \mem_reg_116][17  ( .D(D_17), .E(n6281), .C(wclk), .QN(n3343) );
  DFE1 \mem_reg_116][16  ( .D(D_16), .E(n6281), .C(wclk), .QN(n3344) );
  DFE1 \mem_reg_116][15  ( .D(D_15), .E(n6281), .C(wclk), .QN(n3345) );
  DFE1 \mem_reg_116][14  ( .D(D_14), .E(n6281), .C(wclk), .QN(n3346) );
  DFE1 \mem_reg_116][13  ( .D(D_13), .E(n6281), .C(wclk), .QN(n3347) );
  DFE1 \mem_reg_116][12  ( .D(D_12), .E(n6281), .C(wclk), .QN(n3348) );
  DFE1 \mem_reg_116][11  ( .D(D_11), .E(n6281), .C(wclk), .QN(n3349) );
  DFE1 \mem_reg_116][10  ( .D(D_10), .E(n6281), .C(wclk), .QN(n3350) );
  DFE1 \mem_reg_116][9  ( .D(D_9), .E(n6281), .C(wclk), .QN(n3351) );
  DFE1 \mem_reg_116][8  ( .D(D_8), .E(n6281), .C(wclk), .QN(n3352) );
  DFE1 \mem_reg_116][7  ( .D(D_7), .E(n6281), .C(wclk), .QN(n3353) );
  DFE1 \mem_reg_116][6  ( .D(D_6), .E(n6281), .C(wclk), .QN(n3354) );
  DFE1 \mem_reg_116][5  ( .D(D_5), .E(n6281), .C(wclk), .QN(n3355) );
  DFE1 \mem_reg_116][4  ( .D(D_4), .E(n6281), .C(wclk), .QN(n3356) );
  DFE1 \mem_reg_116][3  ( .D(D_3), .E(n6281), .C(wclk), .QN(n3357) );
  DFE1 \mem_reg_116][2  ( .D(D_2), .E(n6281), .C(wclk), .QN(n3358) );
  DFE1 \mem_reg_116][1  ( .D(D_1), .E(n6281), .C(wclk), .QN(n3359) );
  DFE1 \mem_reg_116][0  ( .D(D_0), .E(n6281), .C(wclk), .QN(n3360) );
  DFE1 \mem_reg_115][23  ( .D(D_23), .E(n6280), .C(wclk), .QN(n3361) );
  DFE1 \mem_reg_115][22  ( .D(D_22), .E(n6280), .C(wclk), .QN(n3362) );
  DFE1 \mem_reg_115][21  ( .D(D_21), .E(n6280), .C(wclk), .QN(n3363) );
  DFE1 \mem_reg_115][20  ( .D(D_20), .E(n6280), .C(wclk), .QN(n3364) );
  DFE1 \mem_reg_115][19  ( .D(D_19), .E(n6280), .C(wclk), .QN(n3365) );
  DFE1 \mem_reg_115][18  ( .D(D_18), .E(n6280), .C(wclk), .QN(n3366) );
  DFE1 \mem_reg_115][17  ( .D(D_17), .E(n6280), .C(wclk), .QN(n3367) );
  DFE1 \mem_reg_115][16  ( .D(D_16), .E(n6280), .C(wclk), .QN(n3368) );
  DFE1 \mem_reg_115][15  ( .D(D_15), .E(n6280), .C(wclk), .QN(n3369) );
  DFE1 \mem_reg_115][14  ( .D(D_14), .E(n6280), .C(wclk), .QN(n3370) );
  DFE1 \mem_reg_115][13  ( .D(D_13), .E(n6280), .C(wclk), .QN(n3371) );
  DFE1 \mem_reg_115][12  ( .D(D_12), .E(n6280), .C(wclk), .QN(n3372) );
  DFE1 \mem_reg_115][11  ( .D(D_11), .E(n6280), .C(wclk), .QN(n3373) );
  DFE1 \mem_reg_115][10  ( .D(D_10), .E(n6280), .C(wclk), .QN(n3374) );
  DFE1 \mem_reg_115][9  ( .D(D_9), .E(n6280), .C(wclk), .QN(n3375) );
  DFE1 \mem_reg_115][8  ( .D(D_8), .E(n6280), .C(wclk), .QN(n3376) );
  DFE1 \mem_reg_115][7  ( .D(D_7), .E(n6280), .C(wclk), .QN(n3377) );
  DFE1 \mem_reg_115][6  ( .D(D_6), .E(n6280), .C(wclk), .QN(n3378) );
  DFE1 \mem_reg_115][5  ( .D(D_5), .E(n6280), .C(wclk), .QN(n3379) );
  DFE1 \mem_reg_115][4  ( .D(D_4), .E(n6280), .C(wclk), .QN(n3380) );
  DFE1 \mem_reg_115][3  ( .D(D_3), .E(n6280), .C(wclk), .QN(n3381) );
  DFE1 \mem_reg_115][2  ( .D(D_2), .E(n6280), .C(wclk), .QN(n3382) );
  DFE1 \mem_reg_115][1  ( .D(D_1), .E(n6280), .C(wclk), .QN(n3383) );
  DFE1 \mem_reg_115][0  ( .D(D_0), .E(n6280), .C(wclk), .QN(n3384) );
  DFE1 \mem_reg_114][23  ( .D(D_23), .E(n6279), .C(wclk), .QN(n3385) );
  DFE1 \mem_reg_114][22  ( .D(D_22), .E(n6279), .C(wclk), .QN(n3386) );
  DFE1 \mem_reg_114][21  ( .D(D_21), .E(n6279), .C(wclk), .QN(n3387) );
  DFE1 \mem_reg_114][20  ( .D(D_20), .E(n6279), .C(wclk), .QN(n3388) );
  DFE1 \mem_reg_114][19  ( .D(D_19), .E(n6279), .C(wclk), .QN(n3389) );
  DFE1 \mem_reg_114][18  ( .D(D_18), .E(n6279), .C(wclk), .QN(n3390) );
  DFE1 \mem_reg_114][17  ( .D(D_17), .E(n6279), .C(wclk), .QN(n3391) );
  DFE1 \mem_reg_114][16  ( .D(D_16), .E(n6279), .C(wclk), .QN(n3392) );
  DFE1 \mem_reg_114][15  ( .D(D_15), .E(n6279), .C(wclk), .QN(n3393) );
  DFE1 \mem_reg_114][14  ( .D(D_14), .E(n6279), .C(wclk), .QN(n3394) );
  DFE1 \mem_reg_114][13  ( .D(D_13), .E(n6279), .C(wclk), .QN(n3395) );
  DFE1 \mem_reg_114][12  ( .D(D_12), .E(n6279), .C(wclk), .QN(n3396) );
  DFE1 \mem_reg_114][11  ( .D(D_11), .E(n6279), .C(wclk), .QN(n3397) );
  DFE1 \mem_reg_114][10  ( .D(D_10), .E(n6279), .C(wclk), .QN(n3398) );
  DFE1 \mem_reg_114][9  ( .D(D_9), .E(n6279), .C(wclk), .QN(n3399) );
  DFE1 \mem_reg_114][8  ( .D(D_8), .E(n6279), .C(wclk), .QN(n3400) );
  DFE1 \mem_reg_114][7  ( .D(D_7), .E(n6279), .C(wclk), .QN(n3401) );
  DFE1 \mem_reg_114][6  ( .D(D_6), .E(n6279), .C(wclk), .QN(n3402) );
  DFE1 \mem_reg_114][5  ( .D(D_5), .E(n6279), .C(wclk), .QN(n3403) );
  DFE1 \mem_reg_114][4  ( .D(D_4), .E(n6279), .C(wclk), .QN(n3404) );
  DFE1 \mem_reg_114][3  ( .D(D_3), .E(n6279), .C(wclk), .QN(n3405) );
  DFE1 \mem_reg_114][2  ( .D(D_2), .E(n6279), .C(wclk), .QN(n3406) );
  DFE1 \mem_reg_114][1  ( .D(D_1), .E(n6279), .C(wclk), .QN(n3407) );
  DFE1 \mem_reg_114][0  ( .D(D_0), .E(n6279), .C(wclk), .QN(n3408) );
  DFE1 \mem_reg_113][23  ( .D(D_23), .E(n6277), .C(wclk), .QN(n3409) );
  DFE1 \mem_reg_113][22  ( .D(D_22), .E(n6277), .C(wclk), .QN(n3410) );
  DFE1 \mem_reg_113][21  ( .D(D_21), .E(n6277), .C(wclk), .QN(n3411) );
  DFE1 \mem_reg_113][20  ( .D(D_20), .E(n6277), .C(wclk), .QN(n3412) );
  DFE1 \mem_reg_113][19  ( .D(D_19), .E(n6277), .C(wclk), .QN(n3413) );
  DFE1 \mem_reg_113][18  ( .D(D_18), .E(n6277), .C(wclk), .QN(n3414) );
  DFE1 \mem_reg_113][17  ( .D(D_17), .E(n6277), .C(wclk), .QN(n3415) );
  DFE1 \mem_reg_113][16  ( .D(D_16), .E(n6277), .C(wclk), .QN(n3416) );
  DFE1 \mem_reg_113][15  ( .D(D_15), .E(n6277), .C(wclk), .QN(n3417) );
  DFE1 \mem_reg_113][14  ( .D(D_14), .E(n6277), .C(wclk), .QN(n3418) );
  DFE1 \mem_reg_113][13  ( .D(D_13), .E(n6277), .C(wclk), .QN(n3419) );
  DFE1 \mem_reg_113][12  ( .D(D_12), .E(n6277), .C(wclk), .QN(n3420) );
  DFE1 \mem_reg_113][11  ( .D(D_11), .E(n6277), .C(wclk), .QN(n3421) );
  DFE1 \mem_reg_113][10  ( .D(D_10), .E(n6277), .C(wclk), .QN(n3422) );
  DFE1 \mem_reg_113][9  ( .D(D_9), .E(n6277), .C(wclk), .QN(n3423) );
  DFE1 \mem_reg_113][8  ( .D(D_8), .E(n6277), .C(wclk), .QN(n3424) );
  DFE1 \mem_reg_113][7  ( .D(D_7), .E(n6277), .C(wclk), .QN(n3425) );
  DFE1 \mem_reg_113][6  ( .D(D_6), .E(n6277), .C(wclk), .QN(n3426) );
  DFE1 \mem_reg_113][5  ( .D(D_5), .E(n6277), .C(wclk), .QN(n3427) );
  DFE1 \mem_reg_113][4  ( .D(D_4), .E(n6277), .C(wclk), .QN(n3428) );
  DFE1 \mem_reg_113][3  ( .D(D_3), .E(n6277), .C(wclk), .QN(n3429) );
  DFE1 \mem_reg_113][2  ( .D(D_2), .E(n6277), .C(wclk), .QN(n3430) );
  DFE1 \mem_reg_113][1  ( .D(D_1), .E(n6277), .C(wclk), .QN(n3431) );
  DFE1 \mem_reg_113][0  ( .D(D_0), .E(n6277), .C(wclk), .QN(n3432) );
  DFE1 \mem_reg_112][23  ( .D(D_23), .E(n6275), .C(wclk), .QN(n3433) );
  DFE1 \mem_reg_112][22  ( .D(D_22), .E(n6275), .C(wclk), .QN(n3434) );
  DFE1 \mem_reg_112][21  ( .D(D_21), .E(n6275), .C(wclk), .QN(n3435) );
  DFE1 \mem_reg_112][20  ( .D(D_20), .E(n6275), .C(wclk), .QN(n3436) );
  DFE1 \mem_reg_112][19  ( .D(D_19), .E(n6275), .C(wclk), .QN(n3437) );
  DFE1 \mem_reg_112][18  ( .D(D_18), .E(n6275), .C(wclk), .QN(n3438) );
  DFE1 \mem_reg_112][17  ( .D(D_17), .E(n6275), .C(wclk), .QN(n3439) );
  DFE1 \mem_reg_112][16  ( .D(D_16), .E(n6275), .C(wclk), .QN(n3440) );
  DFE1 \mem_reg_112][15  ( .D(D_15), .E(n6275), .C(wclk), .QN(n3441) );
  DFE1 \mem_reg_112][14  ( .D(D_14), .E(n6275), .C(wclk), .QN(n3442) );
  DFE1 \mem_reg_112][13  ( .D(D_13), .E(n6275), .C(wclk), .QN(n3443) );
  DFE1 \mem_reg_112][12  ( .D(D_12), .E(n6275), .C(wclk), .QN(n3444) );
  DFE1 \mem_reg_112][11  ( .D(D_11), .E(n6275), .C(wclk), .QN(n3445) );
  DFE1 \mem_reg_112][10  ( .D(D_10), .E(n6275), .C(wclk), .QN(n3446) );
  DFE1 \mem_reg_112][9  ( .D(D_9), .E(n6275), .C(wclk), .QN(n3447) );
  DFE1 \mem_reg_112][8  ( .D(D_8), .E(n6275), .C(wclk), .QN(n3448) );
  DFE1 \mem_reg_112][7  ( .D(D_7), .E(n6275), .C(wclk), .QN(n3449) );
  DFE1 \mem_reg_112][6  ( .D(D_6), .E(n6275), .C(wclk), .QN(n3450) );
  DFE1 \mem_reg_112][5  ( .D(D_5), .E(n6275), .C(wclk), .QN(n3451) );
  DFE1 \mem_reg_112][4  ( .D(D_4), .E(n6275), .C(wclk), .QN(n3452) );
  DFE1 \mem_reg_112][3  ( .D(D_3), .E(n6275), .C(wclk), .QN(n3453) );
  DFE1 \mem_reg_112][2  ( .D(D_2), .E(n6275), .C(wclk), .QN(n3454) );
  DFE1 \mem_reg_112][1  ( .D(D_1), .E(n6275), .C(wclk), .QN(n3455) );
  DFE1 \mem_reg_112][0  ( .D(D_0), .E(n6275), .C(wclk), .QN(n3456) );
  DFE1 \mem_reg_79][23  ( .D(D_23), .E(n6233), .C(wclk), .QN(n4225) );
  DFE1 \mem_reg_79][22  ( .D(D_22), .E(n6233), .C(wclk), .QN(n4226) );
  DFE1 \mem_reg_79][21  ( .D(D_21), .E(n6233), .C(wclk), .QN(n4227) );
  DFE1 \mem_reg_79][20  ( .D(D_20), .E(n6233), .C(wclk), .QN(n4228) );
  DFE1 \mem_reg_79][19  ( .D(D_19), .E(n6233), .C(wclk), .QN(n4229) );
  DFE1 \mem_reg_79][18  ( .D(D_18), .E(n6233), .C(wclk), .QN(n4230) );
  DFE1 \mem_reg_79][17  ( .D(D_17), .E(n6233), .C(wclk), .QN(n4231) );
  DFE1 \mem_reg_79][16  ( .D(D_16), .E(n6233), .C(wclk), .QN(n4232) );
  DFE1 \mem_reg_79][15  ( .D(D_15), .E(n6233), .C(wclk), .QN(n4233) );
  DFE1 \mem_reg_79][14  ( .D(D_14), .E(n6233), .C(wclk), .QN(n4234) );
  DFE1 \mem_reg_79][13  ( .D(D_13), .E(n6233), .C(wclk), .QN(n4235) );
  DFE1 \mem_reg_79][12  ( .D(D_12), .E(n6233), .C(wclk), .QN(n4236) );
  DFE1 \mem_reg_79][11  ( .D(D_11), .E(n6233), .C(wclk), .QN(n4237) );
  DFE1 \mem_reg_79][10  ( .D(D_10), .E(n6233), .C(wclk), .QN(n4238) );
  DFE1 \mem_reg_79][9  ( .D(D_9), .E(n6233), .C(wclk), .QN(n4239) );
  DFE1 \mem_reg_79][8  ( .D(D_8), .E(n6233), .C(wclk), .QN(n4240) );
  DFE1 \mem_reg_79][7  ( .D(D_7), .E(n6233), .C(wclk), .QN(n4241) );
  DFE1 \mem_reg_79][6  ( .D(D_6), .E(n6233), .C(wclk), .QN(n4242) );
  DFE1 \mem_reg_79][5  ( .D(D_5), .E(n6233), .C(wclk), .QN(n4243) );
  DFE1 \mem_reg_79][4  ( .D(D_4), .E(n6233), .C(wclk), .QN(n4244) );
  DFE1 \mem_reg_79][3  ( .D(D_3), .E(n6233), .C(wclk), .QN(n4245) );
  DFE1 \mem_reg_79][2  ( .D(D_2), .E(n6233), .C(wclk), .QN(n4246) );
  DFE1 \mem_reg_79][1  ( .D(D_1), .E(n6233), .C(wclk), .QN(n4247) );
  DFE1 \mem_reg_79][0  ( .D(D_0), .E(n6233), .C(wclk), .QN(n4248) );
  DFE1 \mem_reg_78][23  ( .D(D_23), .E(n6232), .C(wclk), .QN(n4249) );
  DFE1 \mem_reg_78][22  ( .D(D_22), .E(n6232), .C(wclk), .QN(n4250) );
  DFE1 \mem_reg_78][21  ( .D(D_21), .E(n6232), .C(wclk), .QN(n4251) );
  DFE1 \mem_reg_78][20  ( .D(D_20), .E(n6232), .C(wclk), .QN(n4252) );
  DFE1 \mem_reg_78][19  ( .D(D_19), .E(n6232), .C(wclk), .QN(n4253) );
  DFE1 \mem_reg_78][18  ( .D(D_18), .E(n6232), .C(wclk), .QN(n4254) );
  DFE1 \mem_reg_78][17  ( .D(D_17), .E(n6232), .C(wclk), .QN(n4255) );
  DFE1 \mem_reg_78][16  ( .D(D_16), .E(n6232), .C(wclk), .QN(n4256) );
  DFE1 \mem_reg_78][15  ( .D(D_15), .E(n6232), .C(wclk), .QN(n4257) );
  DFE1 \mem_reg_78][14  ( .D(D_14), .E(n6232), .C(wclk), .QN(n4258) );
  DFE1 \mem_reg_78][13  ( .D(D_13), .E(n6232), .C(wclk), .QN(n4259) );
  DFE1 \mem_reg_78][12  ( .D(D_12), .E(n6232), .C(wclk), .QN(n4260) );
  DFE1 \mem_reg_78][11  ( .D(D_11), .E(n6232), .C(wclk), .QN(n4261) );
  DFE1 \mem_reg_78][10  ( .D(D_10), .E(n6232), .C(wclk), .QN(n4262) );
  DFE1 \mem_reg_78][9  ( .D(D_9), .E(n6232), .C(wclk), .QN(n4263) );
  DFE1 \mem_reg_78][8  ( .D(D_8), .E(n6232), .C(wclk), .QN(n4264) );
  DFE1 \mem_reg_78][7  ( .D(D_7), .E(n6232), .C(wclk), .QN(n4265) );
  DFE1 \mem_reg_78][6  ( .D(D_6), .E(n6232), .C(wclk), .QN(n4266) );
  DFE1 \mem_reg_78][5  ( .D(D_5), .E(n6232), .C(wclk), .QN(n4267) );
  DFE1 \mem_reg_78][4  ( .D(D_4), .E(n6232), .C(wclk), .QN(n4268) );
  DFE1 \mem_reg_78][3  ( .D(D_3), .E(n6232), .C(wclk), .QN(n4269) );
  DFE1 \mem_reg_78][2  ( .D(D_2), .E(n6232), .C(wclk), .QN(n4270) );
  DFE1 \mem_reg_78][1  ( .D(D_1), .E(n6232), .C(wclk), .QN(n4271) );
  DFE1 \mem_reg_78][0  ( .D(D_0), .E(n6232), .C(wclk), .QN(n4272) );
  DFE1 \mem_reg_77][23  ( .D(D_23), .E(n6230), .C(wclk), .QN(n4273) );
  DFE1 \mem_reg_77][22  ( .D(D_22), .E(n6230), .C(wclk), .QN(n4274) );
  DFE1 \mem_reg_77][21  ( .D(D_21), .E(n6230), .C(wclk), .QN(n4275) );
  DFE1 \mem_reg_77][20  ( .D(D_20), .E(n6230), .C(wclk), .QN(n4276) );
  DFE1 \mem_reg_77][19  ( .D(D_19), .E(n6230), .C(wclk), .QN(n4277) );
  DFE1 \mem_reg_77][18  ( .D(D_18), .E(n6230), .C(wclk), .QN(n4278) );
  DFE1 \mem_reg_77][17  ( .D(D_17), .E(n6230), .C(wclk), .QN(n4279) );
  DFE1 \mem_reg_77][16  ( .D(D_16), .E(n6230), .C(wclk), .QN(n4280) );
  DFE1 \mem_reg_77][15  ( .D(D_15), .E(n6230), .C(wclk), .QN(n4281) );
  DFE1 \mem_reg_77][14  ( .D(D_14), .E(n6230), .C(wclk), .QN(n4282) );
  DFE1 \mem_reg_77][13  ( .D(D_13), .E(n6230), .C(wclk), .QN(n4283) );
  DFE1 \mem_reg_77][12  ( .D(D_12), .E(n6230), .C(wclk), .QN(n4284) );
  DFE1 \mem_reg_77][11  ( .D(D_11), .E(n6230), .C(wclk), .QN(n4285) );
  DFE1 \mem_reg_77][10  ( .D(D_10), .E(n6230), .C(wclk), .QN(n4286) );
  DFE1 \mem_reg_77][9  ( .D(D_9), .E(n6230), .C(wclk), .QN(n4287) );
  DFE1 \mem_reg_77][8  ( .D(D_8), .E(n6230), .C(wclk), .QN(n4288) );
  DFE1 \mem_reg_77][7  ( .D(D_7), .E(n6230), .C(wclk), .QN(n4289) );
  DFE1 \mem_reg_77][6  ( .D(D_6), .E(n6230), .C(wclk), .QN(n4290) );
  DFE1 \mem_reg_77][5  ( .D(D_5), .E(n6230), .C(wclk), .QN(n4291) );
  DFE1 \mem_reg_77][4  ( .D(D_4), .E(n6230), .C(wclk), .QN(n4292) );
  DFE1 \mem_reg_77][3  ( .D(D_3), .E(n6230), .C(wclk), .QN(n4293) );
  DFE1 \mem_reg_77][2  ( .D(D_2), .E(n6230), .C(wclk), .QN(n4294) );
  DFE1 \mem_reg_77][1  ( .D(D_1), .E(n6230), .C(wclk), .QN(n4295) );
  DFE1 \mem_reg_77][0  ( .D(D_0), .E(n6230), .C(wclk), .QN(n4296) );
  DFE1 \mem_reg_73][23  ( .D(D_23), .E(n6220), .C(wclk), .QN(n4369) );
  DFE1 \mem_reg_73][22  ( .D(D_22), .E(n6220), .C(wclk), .QN(n4370) );
  DFE1 \mem_reg_73][21  ( .D(D_21), .E(n6220), .C(wclk), .QN(n4371) );
  DFE1 \mem_reg_73][20  ( .D(D_20), .E(n6220), .C(wclk), .QN(n4372) );
  DFE1 \mem_reg_73][19  ( .D(D_19), .E(n6220), .C(wclk), .QN(n4373) );
  DFE1 \mem_reg_73][18  ( .D(D_18), .E(n6220), .C(wclk), .QN(n4374) );
  DFE1 \mem_reg_73][17  ( .D(D_17), .E(n6220), .C(wclk), .QN(n4375) );
  DFE1 \mem_reg_73][16  ( .D(D_16), .E(n6220), .C(wclk), .QN(n4376) );
  DFE1 \mem_reg_73][15  ( .D(D_15), .E(n6220), .C(wclk), .QN(n4377) );
  DFE1 \mem_reg_73][14  ( .D(D_14), .E(n6220), .C(wclk), .QN(n4378) );
  DFE1 \mem_reg_73][13  ( .D(D_13), .E(n6220), .C(wclk), .QN(n4379) );
  DFE1 \mem_reg_73][12  ( .D(D_12), .E(n6220), .C(wclk), .QN(n4380) );
  DFE1 \mem_reg_73][11  ( .D(D_11), .E(n6220), .C(wclk), .QN(n4381) );
  DFE1 \mem_reg_73][10  ( .D(D_10), .E(n6220), .C(wclk), .QN(n4382) );
  DFE1 \mem_reg_73][9  ( .D(D_9), .E(n6220), .C(wclk), .QN(n4383) );
  DFE1 \mem_reg_73][8  ( .D(D_8), .E(n6220), .C(wclk), .QN(n4384) );
  DFE1 \mem_reg_73][7  ( .D(D_7), .E(n6220), .C(wclk), .QN(n4385) );
  DFE1 \mem_reg_73][6  ( .D(D_6), .E(n6220), .C(wclk), .QN(n4386) );
  DFE1 \mem_reg_73][5  ( .D(D_5), .E(n6220), .C(wclk), .QN(n4387) );
  DFE1 \mem_reg_73][4  ( .D(D_4), .E(n6220), .C(wclk), .QN(n4388) );
  DFE1 \mem_reg_73][3  ( .D(D_3), .E(n6220), .C(wclk), .QN(n4389) );
  DFE1 \mem_reg_73][2  ( .D(D_2), .E(n6220), .C(wclk), .QN(n4390) );
  DFE1 \mem_reg_73][1  ( .D(D_1), .E(n6220), .C(wclk), .QN(n4391) );
  DFE1 \mem_reg_73][0  ( .D(D_0), .E(n6220), .C(wclk), .QN(n4392) );
  DFE1 \mem_reg_72][23  ( .D(D_23), .E(n6218), .C(wclk), .QN(n4393) );
  DFE1 \mem_reg_72][22  ( .D(D_22), .E(n6218), .C(wclk), .QN(n4394) );
  DFE1 \mem_reg_72][21  ( .D(D_21), .E(n6218), .C(wclk), .QN(n4395) );
  DFE1 \mem_reg_72][20  ( .D(D_20), .E(n6218), .C(wclk), .QN(n4396) );
  DFE1 \mem_reg_72][19  ( .D(D_19), .E(n6218), .C(wclk), .QN(n4397) );
  DFE1 \mem_reg_72][18  ( .D(D_18), .E(n6218), .C(wclk), .QN(n4398) );
  DFE1 \mem_reg_72][17  ( .D(D_17), .E(n6218), .C(wclk), .QN(n4399) );
  DFE1 \mem_reg_72][16  ( .D(D_16), .E(n6218), .C(wclk), .QN(n4400) );
  DFE1 \mem_reg_72][15  ( .D(D_15), .E(n6218), .C(wclk), .QN(n4401) );
  DFE1 \mem_reg_72][14  ( .D(D_14), .E(n6218), .C(wclk), .QN(n4402) );
  DFE1 \mem_reg_72][13  ( .D(D_13), .E(n6218), .C(wclk), .QN(n4403) );
  DFE1 \mem_reg_72][12  ( .D(D_12), .E(n6218), .C(wclk), .QN(n4404) );
  DFE1 \mem_reg_72][11  ( .D(D_11), .E(n6218), .C(wclk), .QN(n4405) );
  DFE1 \mem_reg_72][10  ( .D(D_10), .E(n6218), .C(wclk), .QN(n4406) );
  DFE1 \mem_reg_72][9  ( .D(D_9), .E(n6218), .C(wclk), .QN(n4407) );
  DFE1 \mem_reg_72][8  ( .D(D_8), .E(n6218), .C(wclk), .QN(n4408) );
  DFE1 \mem_reg_72][7  ( .D(D_7), .E(n6218), .C(wclk), .QN(n4409) );
  DFE1 \mem_reg_72][6  ( .D(D_6), .E(n6218), .C(wclk), .QN(n4410) );
  DFE1 \mem_reg_72][5  ( .D(D_5), .E(n6218), .C(wclk), .QN(n4411) );
  DFE1 \mem_reg_72][4  ( .D(D_4), .E(n6218), .C(wclk), .QN(n4412) );
  DFE1 \mem_reg_72][3  ( .D(D_3), .E(n6218), .C(wclk), .QN(n4413) );
  DFE1 \mem_reg_72][2  ( .D(D_2), .E(n6218), .C(wclk), .QN(n4414) );
  DFE1 \mem_reg_72][1  ( .D(D_1), .E(n6218), .C(wclk), .QN(n4415) );
  DFE1 \mem_reg_72][0  ( .D(D_0), .E(n6218), .C(wclk), .QN(n4416) );
  DFE1 \mem_reg_64][23  ( .D(D_23), .E(n6201), .C(wclk), .QN(n4585) );
  DFE1 \mem_reg_64][22  ( .D(D_22), .E(n6201), .C(wclk), .QN(n4586) );
  DFE1 \mem_reg_64][21  ( .D(D_21), .E(n6201), .C(wclk), .QN(n4587) );
  DFE1 \mem_reg_64][20  ( .D(D_20), .E(n6201), .C(wclk), .QN(n4588) );
  DFE1 \mem_reg_64][19  ( .D(D_19), .E(n6201), .C(wclk), .QN(n4589) );
  DFE1 \mem_reg_64][18  ( .D(D_18), .E(n6201), .C(wclk), .QN(n4590) );
  DFE1 \mem_reg_64][17  ( .D(D_17), .E(n6201), .C(wclk), .QN(n4591) );
  DFE1 \mem_reg_64][16  ( .D(D_16), .E(n6201), .C(wclk), .QN(n4592) );
  DFE1 \mem_reg_64][15  ( .D(D_15), .E(n6201), .C(wclk), .QN(n4593) );
  DFE1 \mem_reg_64][14  ( .D(D_14), .E(n6201), .C(wclk), .QN(n4594) );
  DFE1 \mem_reg_64][13  ( .D(D_13), .E(n6201), .C(wclk), .QN(n4595) );
  DFE1 \mem_reg_64][12  ( .D(D_12), .E(n6201), .C(wclk), .QN(n4596) );
  DFE1 \mem_reg_64][11  ( .D(D_11), .E(n6201), .C(wclk), .QN(n4597) );
  DFE1 \mem_reg_64][10  ( .D(D_10), .E(n6201), .C(wclk), .QN(n4598) );
  DFE1 \mem_reg_64][9  ( .D(D_9), .E(n6201), .C(wclk), .QN(n4599) );
  DFE1 \mem_reg_64][8  ( .D(D_8), .E(n6201), .C(wclk), .QN(n4600) );
  DFE1 \mem_reg_64][7  ( .D(D_7), .E(n6201), .C(wclk), .QN(n4601) );
  DFE1 \mem_reg_64][6  ( .D(D_6), .E(n6201), .C(wclk), .QN(n4602) );
  DFE1 \mem_reg_64][5  ( .D(D_5), .E(n6201), .C(wclk), .QN(n4603) );
  DFE1 \mem_reg_64][4  ( .D(D_4), .E(n6201), .C(wclk), .QN(n4604) );
  DFE1 \mem_reg_64][3  ( .D(D_3), .E(n6201), .C(wclk), .QN(n4605) );
  DFE1 \mem_reg_64][2  ( .D(D_2), .E(n6201), .C(wclk), .QN(n4606) );
  DFE1 \mem_reg_64][1  ( .D(D_1), .E(n6201), .C(wclk), .QN(n4607) );
  DFE1 \mem_reg_64][0  ( .D(D_0), .E(n6201), .C(wclk), .QN(n4608) );
  DFE1 \mem_reg_239][23  ( .D(D_23), .E(n6415), .C(wclk), .QN(n385) );
  DFE1 \mem_reg_239][22  ( .D(D_22), .E(n6415), .C(wclk), .QN(n386) );
  DFE1 \mem_reg_239][21  ( .D(D_21), .E(n6415), .C(wclk), .QN(n387) );
  DFE1 \mem_reg_239][20  ( .D(D_20), .E(n6415), .C(wclk), .QN(n388) );
  DFE1 \mem_reg_239][19  ( .D(D_19), .E(n6415), .C(wclk), .QN(n389) );
  DFE1 \mem_reg_239][18  ( .D(D_18), .E(n6415), .C(wclk), .QN(n390) );
  DFE1 \mem_reg_239][17  ( .D(D_17), .E(n6415), .C(wclk), .QN(n391) );
  DFE1 \mem_reg_239][16  ( .D(D_16), .E(n6415), .C(wclk), .QN(n392) );
  DFE1 \mem_reg_239][15  ( .D(D_15), .E(n6415), .C(wclk), .QN(n393) );
  DFE1 \mem_reg_239][14  ( .D(D_14), .E(n6415), .C(wclk), .QN(n394) );
  DFE1 \mem_reg_239][13  ( .D(D_13), .E(n6415), .C(wclk), .QN(n395) );
  DFE1 \mem_reg_239][12  ( .D(D_12), .E(n6415), .C(wclk), .QN(n396) );
  DFE1 \mem_reg_239][11  ( .D(D_11), .E(n6415), .C(wclk), .QN(n397) );
  DFE1 \mem_reg_239][10  ( .D(D_10), .E(n6415), .C(wclk), .QN(n398) );
  DFE1 \mem_reg_239][9  ( .D(D_9), .E(n6415), .C(wclk), .QN(n399) );
  DFE1 \mem_reg_239][8  ( .D(D_8), .E(n6415), .C(wclk), .QN(n400) );
  DFE1 \mem_reg_239][7  ( .D(D_7), .E(n6415), .C(wclk), .QN(n401) );
  DFE1 \mem_reg_239][6  ( .D(D_6), .E(n6415), .C(wclk), .QN(n402) );
  DFE1 \mem_reg_239][5  ( .D(D_5), .E(n6415), .C(wclk), .QN(n403) );
  DFE1 \mem_reg_239][4  ( .D(D_4), .E(n6415), .C(wclk), .QN(n404) );
  DFE1 \mem_reg_239][3  ( .D(D_3), .E(n6415), .C(wclk), .QN(n405) );
  DFE1 \mem_reg_239][2  ( .D(D_2), .E(n6415), .C(wclk), .QN(n406) );
  DFE1 \mem_reg_239][1  ( .D(D_1), .E(n6415), .C(wclk), .QN(n407) );
  DFE1 \mem_reg_239][0  ( .D(D_0), .E(n6415), .C(wclk), .QN(n408) );
  DFE1 \mem_reg_238][23  ( .D(D_23), .E(n6414), .C(wclk), .QN(n409) );
  DFE1 \mem_reg_238][22  ( .D(D_22), .E(n6414), .C(wclk), .QN(n410) );
  DFE1 \mem_reg_238][21  ( .D(D_21), .E(n6414), .C(wclk), .QN(n411) );
  DFE1 \mem_reg_238][20  ( .D(D_20), .E(n6414), .C(wclk), .QN(n412) );
  DFE1 \mem_reg_238][19  ( .D(D_19), .E(n6414), .C(wclk), .QN(n413) );
  DFE1 \mem_reg_238][18  ( .D(D_18), .E(n6414), .C(wclk), .QN(n414) );
  DFE1 \mem_reg_238][17  ( .D(D_17), .E(n6414), .C(wclk), .QN(n415) );
  DFE1 \mem_reg_238][16  ( .D(D_16), .E(n6414), .C(wclk), .QN(n416) );
  DFE1 \mem_reg_238][15  ( .D(D_15), .E(n6414), .C(wclk), .QN(n417) );
  DFE1 \mem_reg_238][14  ( .D(D_14), .E(n6414), .C(wclk), .QN(n418) );
  DFE1 \mem_reg_238][13  ( .D(D_13), .E(n6414), .C(wclk), .QN(n419) );
  DFE1 \mem_reg_238][12  ( .D(D_12), .E(n6414), .C(wclk), .QN(n420) );
  DFE1 \mem_reg_238][11  ( .D(D_11), .E(n6414), .C(wclk), .QN(n421) );
  DFE1 \mem_reg_238][10  ( .D(D_10), .E(n6414), .C(wclk), .QN(n422) );
  DFE1 \mem_reg_238][9  ( .D(D_9), .E(n6414), .C(wclk), .QN(n423) );
  DFE1 \mem_reg_238][8  ( .D(D_8), .E(n6414), .C(wclk), .QN(n424) );
  DFE1 \mem_reg_238][7  ( .D(D_7), .E(n6414), .C(wclk), .QN(n425) );
  DFE1 \mem_reg_238][6  ( .D(D_6), .E(n6414), .C(wclk), .QN(n426) );
  DFE1 \mem_reg_238][5  ( .D(D_5), .E(n6414), .C(wclk), .QN(n427) );
  DFE1 \mem_reg_238][4  ( .D(D_4), .E(n6414), .C(wclk), .QN(n428) );
  DFE1 \mem_reg_238][3  ( .D(D_3), .E(n6414), .C(wclk), .QN(n429) );
  DFE1 \mem_reg_238][2  ( .D(D_2), .E(n6414), .C(wclk), .QN(n430) );
  DFE1 \mem_reg_238][1  ( .D(D_1), .E(n6414), .C(wclk), .QN(n431) );
  DFE1 \mem_reg_238][0  ( .D(D_0), .E(n6414), .C(wclk), .QN(n432) );
  DFE1 \mem_reg_237][23  ( .D(D_23), .E(n6413), .C(wclk), .QN(n433) );
  DFE1 \mem_reg_237][22  ( .D(D_22), .E(n6413), .C(wclk), .QN(n434) );
  DFE1 \mem_reg_237][21  ( .D(D_21), .E(n6413), .C(wclk), .QN(n435) );
  DFE1 \mem_reg_237][20  ( .D(D_20), .E(n6413), .C(wclk), .QN(n436) );
  DFE1 \mem_reg_237][19  ( .D(D_19), .E(n6413), .C(wclk), .QN(n437) );
  DFE1 \mem_reg_237][18  ( .D(D_18), .E(n6413), .C(wclk), .QN(n438) );
  DFE1 \mem_reg_237][17  ( .D(D_17), .E(n6413), .C(wclk), .QN(n439) );
  DFE1 \mem_reg_237][16  ( .D(D_16), .E(n6413), .C(wclk), .QN(n440) );
  DFE1 \mem_reg_237][15  ( .D(D_15), .E(n6413), .C(wclk), .QN(n441) );
  DFE1 \mem_reg_237][14  ( .D(D_14), .E(n6413), .C(wclk), .QN(n442) );
  DFE1 \mem_reg_237][13  ( .D(D_13), .E(n6413), .C(wclk), .QN(n443) );
  DFE1 \mem_reg_237][12  ( .D(D_12), .E(n6413), .C(wclk), .QN(n444) );
  DFE1 \mem_reg_237][11  ( .D(D_11), .E(n6413), .C(wclk), .QN(n445) );
  DFE1 \mem_reg_237][10  ( .D(D_10), .E(n6413), .C(wclk), .QN(n446) );
  DFE1 \mem_reg_237][9  ( .D(D_9), .E(n6413), .C(wclk), .QN(n447) );
  DFE1 \mem_reg_237][8  ( .D(D_8), .E(n6413), .C(wclk), .QN(n448) );
  DFE1 \mem_reg_237][7  ( .D(D_7), .E(n6413), .C(wclk), .QN(n449) );
  DFE1 \mem_reg_237][6  ( .D(D_6), .E(n6413), .C(wclk), .QN(n450) );
  DFE1 \mem_reg_237][5  ( .D(D_5), .E(n6413), .C(wclk), .QN(n451) );
  DFE1 \mem_reg_237][4  ( .D(D_4), .E(n6413), .C(wclk), .QN(n452) );
  DFE1 \mem_reg_237][3  ( .D(D_3), .E(n6413), .C(wclk), .QN(n453) );
  DFE1 \mem_reg_237][2  ( .D(D_2), .E(n6413), .C(wclk), .QN(n454) );
  DFE1 \mem_reg_237][1  ( .D(D_1), .E(n6413), .C(wclk), .QN(n455) );
  DFE1 \mem_reg_237][0  ( .D(D_0), .E(n6413), .C(wclk), .QN(n456) );
  DFE1 \mem_reg_236][23  ( .D(D_23), .E(n6412), .C(wclk), .QN(n457) );
  DFE1 \mem_reg_236][22  ( .D(D_22), .E(n6412), .C(wclk), .QN(n458) );
  DFE1 \mem_reg_236][21  ( .D(D_21), .E(n6412), .C(wclk), .QN(n459) );
  DFE1 \mem_reg_236][20  ( .D(D_20), .E(n6412), .C(wclk), .QN(n460) );
  DFE1 \mem_reg_236][19  ( .D(D_19), .E(n6412), .C(wclk), .QN(n461) );
  DFE1 \mem_reg_236][18  ( .D(D_18), .E(n6412), .C(wclk), .QN(n462) );
  DFE1 \mem_reg_236][17  ( .D(D_17), .E(n6412), .C(wclk), .QN(n463) );
  DFE1 \mem_reg_236][16  ( .D(D_16), .E(n6412), .C(wclk), .QN(n464) );
  DFE1 \mem_reg_236][15  ( .D(D_15), .E(n6412), .C(wclk), .QN(n465) );
  DFE1 \mem_reg_236][14  ( .D(D_14), .E(n6412), .C(wclk), .QN(n466) );
  DFE1 \mem_reg_236][13  ( .D(D_13), .E(n6412), .C(wclk), .QN(n467) );
  DFE1 \mem_reg_236][12  ( .D(D_12), .E(n6412), .C(wclk), .QN(n468) );
  DFE1 \mem_reg_236][11  ( .D(D_11), .E(n6412), .C(wclk), .QN(n469) );
  DFE1 \mem_reg_236][10  ( .D(D_10), .E(n6412), .C(wclk), .QN(n470) );
  DFE1 \mem_reg_236][9  ( .D(D_9), .E(n6412), .C(wclk), .QN(n471) );
  DFE1 \mem_reg_236][8  ( .D(D_8), .E(n6412), .C(wclk), .QN(n472) );
  DFE1 \mem_reg_236][7  ( .D(D_7), .E(n6412), .C(wclk), .QN(n473) );
  DFE1 \mem_reg_236][6  ( .D(D_6), .E(n6412), .C(wclk), .QN(n474) );
  DFE1 \mem_reg_236][5  ( .D(D_5), .E(n6412), .C(wclk), .QN(n475) );
  DFE1 \mem_reg_236][4  ( .D(D_4), .E(n6412), .C(wclk), .QN(n476) );
  DFE1 \mem_reg_236][3  ( .D(D_3), .E(n6412), .C(wclk), .QN(n477) );
  DFE1 \mem_reg_236][2  ( .D(D_2), .E(n6412), .C(wclk), .QN(n478) );
  DFE1 \mem_reg_236][1  ( .D(D_1), .E(n6412), .C(wclk), .QN(n479) );
  DFE1 \mem_reg_236][0  ( .D(D_0), .E(n6412), .C(wclk), .QN(n480) );
  DFE1 \mem_reg_235][23  ( .D(D_23), .E(n6411), .C(wclk), .QN(n481) );
  DFE1 \mem_reg_235][22  ( .D(D_22), .E(n6411), .C(wclk), .QN(n482) );
  DFE1 \mem_reg_235][21  ( .D(D_21), .E(n6411), .C(wclk), .QN(n483) );
  DFE1 \mem_reg_235][20  ( .D(D_20), .E(n6411), .C(wclk), .QN(n484) );
  DFE1 \mem_reg_235][19  ( .D(D_19), .E(n6411), .C(wclk), .QN(n485) );
  DFE1 \mem_reg_235][18  ( .D(D_18), .E(n6411), .C(wclk), .QN(n486) );
  DFE1 \mem_reg_235][17  ( .D(D_17), .E(n6411), .C(wclk), .QN(n487) );
  DFE1 \mem_reg_235][16  ( .D(D_16), .E(n6411), .C(wclk), .QN(n488) );
  DFE1 \mem_reg_235][15  ( .D(D_15), .E(n6411), .C(wclk), .QN(n489) );
  DFE1 \mem_reg_235][14  ( .D(D_14), .E(n6411), .C(wclk), .QN(n490) );
  DFE1 \mem_reg_235][13  ( .D(D_13), .E(n6411), .C(wclk), .QN(n491) );
  DFE1 \mem_reg_235][12  ( .D(D_12), .E(n6411), .C(wclk), .QN(n492) );
  DFE1 \mem_reg_235][11  ( .D(D_11), .E(n6411), .C(wclk), .QN(n493) );
  DFE1 \mem_reg_235][10  ( .D(D_10), .E(n6411), .C(wclk), .QN(n494) );
  DFE1 \mem_reg_235][9  ( .D(D_9), .E(n6411), .C(wclk), .QN(n495) );
  DFE1 \mem_reg_235][8  ( .D(D_8), .E(n6411), .C(wclk), .QN(n496) );
  DFE1 \mem_reg_235][7  ( .D(D_7), .E(n6411), .C(wclk), .QN(n497) );
  DFE1 \mem_reg_235][6  ( .D(D_6), .E(n6411), .C(wclk), .QN(n498) );
  DFE1 \mem_reg_235][5  ( .D(D_5), .E(n6411), .C(wclk), .QN(n499) );
  DFE1 \mem_reg_235][4  ( .D(D_4), .E(n6411), .C(wclk), .QN(n500) );
  DFE1 \mem_reg_235][3  ( .D(D_3), .E(n6411), .C(wclk), .QN(n501) );
  DFE1 \mem_reg_235][2  ( .D(D_2), .E(n6411), .C(wclk), .QN(n502) );
  DFE1 \mem_reg_235][1  ( .D(D_1), .E(n6411), .C(wclk), .QN(n503) );
  DFE1 \mem_reg_235][0  ( .D(D_0), .E(n6411), .C(wclk), .QN(n504) );
  DFE1 \mem_reg_234][23  ( .D(D_23), .E(n6410), .C(wclk), .QN(n505) );
  DFE1 \mem_reg_234][22  ( .D(D_22), .E(n6410), .C(wclk), .QN(n506) );
  DFE1 \mem_reg_234][21  ( .D(D_21), .E(n6410), .C(wclk), .QN(n507) );
  DFE1 \mem_reg_234][20  ( .D(D_20), .E(n6410), .C(wclk), .QN(n508) );
  DFE1 \mem_reg_234][19  ( .D(D_19), .E(n6410), .C(wclk), .QN(n509) );
  DFE1 \mem_reg_234][18  ( .D(D_18), .E(n6410), .C(wclk), .QN(n510) );
  DFE1 \mem_reg_234][17  ( .D(D_17), .E(n6410), .C(wclk), .QN(n511) );
  DFE1 \mem_reg_234][16  ( .D(D_16), .E(n6410), .C(wclk), .QN(n512) );
  DFE1 \mem_reg_234][15  ( .D(D_15), .E(n6410), .C(wclk), .QN(n513) );
  DFE1 \mem_reg_234][14  ( .D(D_14), .E(n6410), .C(wclk), .QN(n514) );
  DFE1 \mem_reg_234][13  ( .D(D_13), .E(n6410), .C(wclk), .QN(n515) );
  DFE1 \mem_reg_234][12  ( .D(D_12), .E(n6410), .C(wclk), .QN(n516) );
  DFE1 \mem_reg_234][11  ( .D(D_11), .E(n6410), .C(wclk), .QN(n517) );
  DFE1 \mem_reg_234][10  ( .D(D_10), .E(n6410), .C(wclk), .QN(n518) );
  DFE1 \mem_reg_234][9  ( .D(D_9), .E(n6410), .C(wclk), .QN(n519) );
  DFE1 \mem_reg_234][8  ( .D(D_8), .E(n6410), .C(wclk), .QN(n520) );
  DFE1 \mem_reg_234][7  ( .D(D_7), .E(n6410), .C(wclk), .QN(n521) );
  DFE1 \mem_reg_234][6  ( .D(D_6), .E(n6410), .C(wclk), .QN(n522) );
  DFE1 \mem_reg_234][5  ( .D(D_5), .E(n6410), .C(wclk), .QN(n523) );
  DFE1 \mem_reg_234][4  ( .D(D_4), .E(n6410), .C(wclk), .QN(n524) );
  DFE1 \mem_reg_234][3  ( .D(D_3), .E(n6410), .C(wclk), .QN(n525) );
  DFE1 \mem_reg_234][2  ( .D(D_2), .E(n6410), .C(wclk), .QN(n526) );
  DFE1 \mem_reg_234][1  ( .D(D_1), .E(n6410), .C(wclk), .QN(n527) );
  DFE1 \mem_reg_234][0  ( .D(D_0), .E(n6410), .C(wclk), .QN(n528) );
  DFE1 \mem_reg_233][23  ( .D(D_23), .E(n6409), .C(wclk), .QN(n529) );
  DFE1 \mem_reg_233][22  ( .D(D_22), .E(n6409), .C(wclk), .QN(n530) );
  DFE1 \mem_reg_233][21  ( .D(D_21), .E(n6409), .C(wclk), .QN(n531) );
  DFE1 \mem_reg_233][20  ( .D(D_20), .E(n6409), .C(wclk), .QN(n532) );
  DFE1 \mem_reg_233][19  ( .D(D_19), .E(n6409), .C(wclk), .QN(n533) );
  DFE1 \mem_reg_233][18  ( .D(D_18), .E(n6409), .C(wclk), .QN(n534) );
  DFE1 \mem_reg_233][17  ( .D(D_17), .E(n6409), .C(wclk), .QN(n535) );
  DFE1 \mem_reg_233][16  ( .D(D_16), .E(n6409), .C(wclk), .QN(n536) );
  DFE1 \mem_reg_233][15  ( .D(D_15), .E(n6409), .C(wclk), .QN(n537) );
  DFE1 \mem_reg_233][14  ( .D(D_14), .E(n6409), .C(wclk), .QN(n538) );
  DFE1 \mem_reg_233][13  ( .D(D_13), .E(n6409), .C(wclk), .QN(n539) );
  DFE1 \mem_reg_233][12  ( .D(D_12), .E(n6409), .C(wclk), .QN(n540) );
  DFE1 \mem_reg_233][11  ( .D(D_11), .E(n6409), .C(wclk), .QN(n541) );
  DFE1 \mem_reg_233][10  ( .D(D_10), .E(n6409), .C(wclk), .QN(n542) );
  DFE1 \mem_reg_233][9  ( .D(D_9), .E(n6409), .C(wclk), .QN(n543) );
  DFE1 \mem_reg_233][8  ( .D(D_8), .E(n6409), .C(wclk), .QN(n544) );
  DFE1 \mem_reg_233][7  ( .D(D_7), .E(n6409), .C(wclk), .QN(n545) );
  DFE1 \mem_reg_233][6  ( .D(D_6), .E(n6409), .C(wclk), .QN(n546) );
  DFE1 \mem_reg_233][5  ( .D(D_5), .E(n6409), .C(wclk), .QN(n547) );
  DFE1 \mem_reg_233][4  ( .D(D_4), .E(n6409), .C(wclk), .QN(n548) );
  DFE1 \mem_reg_233][3  ( .D(D_3), .E(n6409), .C(wclk), .QN(n549) );
  DFE1 \mem_reg_233][2  ( .D(D_2), .E(n6409), .C(wclk), .QN(n550) );
  DFE1 \mem_reg_233][1  ( .D(D_1), .E(n6409), .C(wclk), .QN(n551) );
  DFE1 \mem_reg_233][0  ( .D(D_0), .E(n6409), .C(wclk), .QN(n552) );
  DFE1 \mem_reg_232][23  ( .D(D_23), .E(n6408), .C(wclk), .QN(n553) );
  DFE1 \mem_reg_232][22  ( .D(D_22), .E(n6408), .C(wclk), .QN(n554) );
  DFE1 \mem_reg_232][21  ( .D(D_21), .E(n6408), .C(wclk), .QN(n555) );
  DFE1 \mem_reg_232][20  ( .D(D_20), .E(n6408), .C(wclk), .QN(n556) );
  DFE1 \mem_reg_232][19  ( .D(D_19), .E(n6408), .C(wclk), .QN(n557) );
  DFE1 \mem_reg_232][18  ( .D(D_18), .E(n6408), .C(wclk), .QN(n558) );
  DFE1 \mem_reg_232][17  ( .D(D_17), .E(n6408), .C(wclk), .QN(n559) );
  DFE1 \mem_reg_232][16  ( .D(D_16), .E(n6408), .C(wclk), .QN(n560) );
  DFE1 \mem_reg_232][15  ( .D(D_15), .E(n6408), .C(wclk), .QN(n561) );
  DFE1 \mem_reg_232][14  ( .D(D_14), .E(n6408), .C(wclk), .QN(n562) );
  DFE1 \mem_reg_232][13  ( .D(D_13), .E(n6408), .C(wclk), .QN(n563) );
  DFE1 \mem_reg_232][12  ( .D(D_12), .E(n6408), .C(wclk), .QN(n564) );
  DFE1 \mem_reg_232][11  ( .D(D_11), .E(n6408), .C(wclk), .QN(n565) );
  DFE1 \mem_reg_232][10  ( .D(D_10), .E(n6408), .C(wclk), .QN(n566) );
  DFE1 \mem_reg_232][9  ( .D(D_9), .E(n6408), .C(wclk), .QN(n567) );
  DFE1 \mem_reg_232][8  ( .D(D_8), .E(n6408), .C(wclk), .QN(n568) );
  DFE1 \mem_reg_232][7  ( .D(D_7), .E(n6408), .C(wclk), .QN(n569) );
  DFE1 \mem_reg_232][6  ( .D(D_6), .E(n6408), .C(wclk), .QN(n570) );
  DFE1 \mem_reg_232][5  ( .D(D_5), .E(n6408), .C(wclk), .QN(n571) );
  DFE1 \mem_reg_232][4  ( .D(D_4), .E(n6408), .C(wclk), .QN(n572) );
  DFE1 \mem_reg_232][3  ( .D(D_3), .E(n6408), .C(wclk), .QN(n573) );
  DFE1 \mem_reg_232][2  ( .D(D_2), .E(n6408), .C(wclk), .QN(n574) );
  DFE1 \mem_reg_232][1  ( .D(D_1), .E(n6408), .C(wclk), .QN(n575) );
  DFE1 \mem_reg_232][0  ( .D(D_0), .E(n6408), .C(wclk), .QN(n576) );
  DFE1 \mem_reg_231][23  ( .D(D_23), .E(n6407), .C(wclk), .QN(n577) );
  DFE1 \mem_reg_231][22  ( .D(D_22), .E(n6407), .C(wclk), .QN(n578) );
  DFE1 \mem_reg_231][21  ( .D(D_21), .E(n6407), .C(wclk), .QN(n579) );
  DFE1 \mem_reg_231][20  ( .D(D_20), .E(n6407), .C(wclk), .QN(n580) );
  DFE1 \mem_reg_231][19  ( .D(D_19), .E(n6407), .C(wclk), .QN(n581) );
  DFE1 \mem_reg_231][18  ( .D(D_18), .E(n6407), .C(wclk), .QN(n582) );
  DFE1 \mem_reg_231][17  ( .D(D_17), .E(n6407), .C(wclk), .QN(n583) );
  DFE1 \mem_reg_231][16  ( .D(D_16), .E(n6407), .C(wclk), .QN(n584) );
  DFE1 \mem_reg_231][15  ( .D(D_15), .E(n6407), .C(wclk), .QN(n585) );
  DFE1 \mem_reg_231][14  ( .D(D_14), .E(n6407), .C(wclk), .QN(n586) );
  DFE1 \mem_reg_231][13  ( .D(D_13), .E(n6407), .C(wclk), .QN(n587) );
  DFE1 \mem_reg_231][12  ( .D(D_12), .E(n6407), .C(wclk), .QN(n588) );
  DFE1 \mem_reg_231][11  ( .D(D_11), .E(n6407), .C(wclk), .QN(n589) );
  DFE1 \mem_reg_231][10  ( .D(D_10), .E(n6407), .C(wclk), .QN(n590) );
  DFE1 \mem_reg_231][9  ( .D(D_9), .E(n6407), .C(wclk), .QN(n591) );
  DFE1 \mem_reg_231][8  ( .D(D_8), .E(n6407), .C(wclk), .QN(n592) );
  DFE1 \mem_reg_231][7  ( .D(D_7), .E(n6407), .C(wclk), .QN(n593) );
  DFE1 \mem_reg_231][6  ( .D(D_6), .E(n6407), .C(wclk), .QN(n594) );
  DFE1 \mem_reg_231][5  ( .D(D_5), .E(n6407), .C(wclk), .QN(n595) );
  DFE1 \mem_reg_231][4  ( .D(D_4), .E(n6407), .C(wclk), .QN(n596) );
  DFE1 \mem_reg_231][3  ( .D(D_3), .E(n6407), .C(wclk), .QN(n597) );
  DFE1 \mem_reg_231][2  ( .D(D_2), .E(n6407), .C(wclk), .QN(n598) );
  DFE1 \mem_reg_231][1  ( .D(D_1), .E(n6407), .C(wclk), .QN(n599) );
  DFE1 \mem_reg_231][0  ( .D(D_0), .E(n6407), .C(wclk), .QN(n600) );
  DFE1 \mem_reg_230][23  ( .D(D_23), .E(n6406), .C(wclk), .QN(n601) );
  DFE1 \mem_reg_230][22  ( .D(D_22), .E(n6406), .C(wclk), .QN(n602) );
  DFE1 \mem_reg_230][21  ( .D(D_21), .E(n6406), .C(wclk), .QN(n603) );
  DFE1 \mem_reg_230][20  ( .D(D_20), .E(n6406), .C(wclk), .QN(n604) );
  DFE1 \mem_reg_230][19  ( .D(D_19), .E(n6406), .C(wclk), .QN(n605) );
  DFE1 \mem_reg_230][18  ( .D(D_18), .E(n6406), .C(wclk), .QN(n606) );
  DFE1 \mem_reg_230][17  ( .D(D_17), .E(n6406), .C(wclk), .QN(n607) );
  DFE1 \mem_reg_230][16  ( .D(D_16), .E(n6406), .C(wclk), .QN(n608) );
  DFE1 \mem_reg_230][15  ( .D(D_15), .E(n6406), .C(wclk), .QN(n609) );
  DFE1 \mem_reg_230][14  ( .D(D_14), .E(n6406), .C(wclk), .QN(n610) );
  DFE1 \mem_reg_230][13  ( .D(D_13), .E(n6406), .C(wclk), .QN(n611) );
  DFE1 \mem_reg_230][12  ( .D(D_12), .E(n6406), .C(wclk), .QN(n612) );
  DFE1 \mem_reg_230][11  ( .D(D_11), .E(n6406), .C(wclk), .QN(n613) );
  DFE1 \mem_reg_230][10  ( .D(D_10), .E(n6406), .C(wclk), .QN(n614) );
  DFE1 \mem_reg_230][9  ( .D(D_9), .E(n6406), .C(wclk), .QN(n615) );
  DFE1 \mem_reg_230][8  ( .D(D_8), .E(n6406), .C(wclk), .QN(n616) );
  DFE1 \mem_reg_230][7  ( .D(D_7), .E(n6406), .C(wclk), .QN(n617) );
  DFE1 \mem_reg_230][6  ( .D(D_6), .E(n6406), .C(wclk), .QN(n618) );
  DFE1 \mem_reg_230][5  ( .D(D_5), .E(n6406), .C(wclk), .QN(n619) );
  DFE1 \mem_reg_230][4  ( .D(D_4), .E(n6406), .C(wclk), .QN(n620) );
  DFE1 \mem_reg_230][3  ( .D(D_3), .E(n6406), .C(wclk), .QN(n621) );
  DFE1 \mem_reg_230][2  ( .D(D_2), .E(n6406), .C(wclk), .QN(n622) );
  DFE1 \mem_reg_230][1  ( .D(D_1), .E(n6406), .C(wclk), .QN(n623) );
  DFE1 \mem_reg_230][0  ( .D(D_0), .E(n6406), .C(wclk), .QN(n624) );
  DFE1 \mem_reg_229][23  ( .D(D_23), .E(n6405), .C(wclk), .QN(n625) );
  DFE1 \mem_reg_229][22  ( .D(D_22), .E(n6405), .C(wclk), .QN(n626) );
  DFE1 \mem_reg_229][21  ( .D(D_21), .E(n6405), .C(wclk), .QN(n627) );
  DFE1 \mem_reg_229][20  ( .D(D_20), .E(n6405), .C(wclk), .QN(n628) );
  DFE1 \mem_reg_229][19  ( .D(D_19), .E(n6405), .C(wclk), .QN(n629) );
  DFE1 \mem_reg_229][18  ( .D(D_18), .E(n6405), .C(wclk), .QN(n630) );
  DFE1 \mem_reg_229][17  ( .D(D_17), .E(n6405), .C(wclk), .QN(n631) );
  DFE1 \mem_reg_229][16  ( .D(D_16), .E(n6405), .C(wclk), .QN(n632) );
  DFE1 \mem_reg_229][15  ( .D(D_15), .E(n6405), .C(wclk), .QN(n633) );
  DFE1 \mem_reg_229][14  ( .D(D_14), .E(n6405), .C(wclk), .QN(n634) );
  DFE1 \mem_reg_229][13  ( .D(D_13), .E(n6405), .C(wclk), .QN(n635) );
  DFE1 \mem_reg_229][12  ( .D(D_12), .E(n6405), .C(wclk), .QN(n636) );
  DFE1 \mem_reg_229][11  ( .D(D_11), .E(n6405), .C(wclk), .QN(n637) );
  DFE1 \mem_reg_229][10  ( .D(D_10), .E(n6405), .C(wclk), .QN(n638) );
  DFE1 \mem_reg_229][9  ( .D(D_9), .E(n6405), .C(wclk), .QN(n639) );
  DFE1 \mem_reg_229][8  ( .D(D_8), .E(n6405), .C(wclk), .QN(n640) );
  DFE1 \mem_reg_229][7  ( .D(D_7), .E(n6405), .C(wclk), .QN(n641) );
  DFE1 \mem_reg_229][6  ( .D(D_6), .E(n6405), .C(wclk), .QN(n642) );
  DFE1 \mem_reg_229][5  ( .D(D_5), .E(n6405), .C(wclk), .QN(n643) );
  DFE1 \mem_reg_229][4  ( .D(D_4), .E(n6405), .C(wclk), .QN(n644) );
  DFE1 \mem_reg_229][3  ( .D(D_3), .E(n6405), .C(wclk), .QN(n645) );
  DFE1 \mem_reg_229][2  ( .D(D_2), .E(n6405), .C(wclk), .QN(n646) );
  DFE1 \mem_reg_229][1  ( .D(D_1), .E(n6405), .C(wclk), .QN(n647) );
  DFE1 \mem_reg_229][0  ( .D(D_0), .E(n6405), .C(wclk), .QN(n648) );
  DFE1 \mem_reg_228][23  ( .D(D_23), .E(n6404), .C(wclk), .QN(n649) );
  DFE1 \mem_reg_228][22  ( .D(D_22), .E(n6404), .C(wclk), .QN(n650) );
  DFE1 \mem_reg_228][21  ( .D(D_21), .E(n6404), .C(wclk), .QN(n651) );
  DFE1 \mem_reg_228][20  ( .D(D_20), .E(n6404), .C(wclk), .QN(n652) );
  DFE1 \mem_reg_228][19  ( .D(D_19), .E(n6404), .C(wclk), .QN(n653) );
  DFE1 \mem_reg_228][18  ( .D(D_18), .E(n6404), .C(wclk), .QN(n654) );
  DFE1 \mem_reg_228][17  ( .D(D_17), .E(n6404), .C(wclk), .QN(n655) );
  DFE1 \mem_reg_228][16  ( .D(D_16), .E(n6404), .C(wclk), .QN(n656) );
  DFE1 \mem_reg_228][15  ( .D(D_15), .E(n6404), .C(wclk), .QN(n657) );
  DFE1 \mem_reg_228][14  ( .D(D_14), .E(n6404), .C(wclk), .QN(n658) );
  DFE1 \mem_reg_228][13  ( .D(D_13), .E(n6404), .C(wclk), .QN(n659) );
  DFE1 \mem_reg_228][12  ( .D(D_12), .E(n6404), .C(wclk), .QN(n660) );
  DFE1 \mem_reg_228][11  ( .D(D_11), .E(n6404), .C(wclk), .QN(n661) );
  DFE1 \mem_reg_228][10  ( .D(D_10), .E(n6404), .C(wclk), .QN(n662) );
  DFE1 \mem_reg_228][9  ( .D(D_9), .E(n6404), .C(wclk), .QN(n663) );
  DFE1 \mem_reg_228][8  ( .D(D_8), .E(n6404), .C(wclk), .QN(n664) );
  DFE1 \mem_reg_228][7  ( .D(D_7), .E(n6404), .C(wclk), .QN(n665) );
  DFE1 \mem_reg_228][6  ( .D(D_6), .E(n6404), .C(wclk), .QN(n666) );
  DFE1 \mem_reg_228][5  ( .D(D_5), .E(n6404), .C(wclk), .QN(n667) );
  DFE1 \mem_reg_228][4  ( .D(D_4), .E(n6404), .C(wclk), .QN(n668) );
  DFE1 \mem_reg_228][3  ( .D(D_3), .E(n6404), .C(wclk), .QN(n669) );
  DFE1 \mem_reg_228][2  ( .D(D_2), .E(n6404), .C(wclk), .QN(n670) );
  DFE1 \mem_reg_228][1  ( .D(D_1), .E(n6404), .C(wclk), .QN(n671) );
  DFE1 \mem_reg_228][0  ( .D(D_0), .E(n6404), .C(wclk), .QN(n672) );
  DFE1 \mem_reg_227][23  ( .D(D_23), .E(n6403), .C(wclk), .QN(n673) );
  DFE1 \mem_reg_227][22  ( .D(D_22), .E(n6403), .C(wclk), .QN(n674) );
  DFE1 \mem_reg_227][21  ( .D(D_21), .E(n6403), .C(wclk), .QN(n675) );
  DFE1 \mem_reg_227][20  ( .D(D_20), .E(n6403), .C(wclk), .QN(n676) );
  DFE1 \mem_reg_227][19  ( .D(D_19), .E(n6403), .C(wclk), .QN(n677) );
  DFE1 \mem_reg_227][18  ( .D(D_18), .E(n6403), .C(wclk), .QN(n678) );
  DFE1 \mem_reg_227][17  ( .D(D_17), .E(n6403), .C(wclk), .QN(n679) );
  DFE1 \mem_reg_227][16  ( .D(D_16), .E(n6403), .C(wclk), .QN(n680) );
  DFE1 \mem_reg_227][15  ( .D(D_15), .E(n6403), .C(wclk), .QN(n681) );
  DFE1 \mem_reg_227][14  ( .D(D_14), .E(n6403), .C(wclk), .QN(n682) );
  DFE1 \mem_reg_227][13  ( .D(D_13), .E(n6403), .C(wclk), .QN(n683) );
  DFE1 \mem_reg_227][12  ( .D(D_12), .E(n6403), .C(wclk), .QN(n684) );
  DFE1 \mem_reg_227][11  ( .D(D_11), .E(n6403), .C(wclk), .QN(n685) );
  DFE1 \mem_reg_227][10  ( .D(D_10), .E(n6403), .C(wclk), .QN(n686) );
  DFE1 \mem_reg_227][9  ( .D(D_9), .E(n6403), .C(wclk), .QN(n687) );
  DFE1 \mem_reg_227][8  ( .D(D_8), .E(n6403), .C(wclk), .QN(n688) );
  DFE1 \mem_reg_227][7  ( .D(D_7), .E(n6403), .C(wclk), .QN(n689) );
  DFE1 \mem_reg_227][6  ( .D(D_6), .E(n6403), .C(wclk), .QN(n690) );
  DFE1 \mem_reg_227][5  ( .D(D_5), .E(n6403), .C(wclk), .QN(n691) );
  DFE1 \mem_reg_227][4  ( .D(D_4), .E(n6403), .C(wclk), .QN(n692) );
  DFE1 \mem_reg_227][3  ( .D(D_3), .E(n6403), .C(wclk), .QN(n693) );
  DFE1 \mem_reg_227][2  ( .D(D_2), .E(n6403), .C(wclk), .QN(n694) );
  DFE1 \mem_reg_227][1  ( .D(D_1), .E(n6403), .C(wclk), .QN(n695) );
  DFE1 \mem_reg_227][0  ( .D(D_0), .E(n6403), .C(wclk), .QN(n696) );
  DFE1 \mem_reg_226][23  ( .D(D_23), .E(n6402), .C(wclk), .QN(n697) );
  DFE1 \mem_reg_226][22  ( .D(D_22), .E(n6402), .C(wclk), .QN(n698) );
  DFE1 \mem_reg_226][21  ( .D(D_21), .E(n6402), .C(wclk), .QN(n699) );
  DFE1 \mem_reg_226][20  ( .D(D_20), .E(n6402), .C(wclk), .QN(n700) );
  DFE1 \mem_reg_226][19  ( .D(D_19), .E(n6402), .C(wclk), .QN(n701) );
  DFE1 \mem_reg_226][18  ( .D(D_18), .E(n6402), .C(wclk), .QN(n702) );
  DFE1 \mem_reg_226][17  ( .D(D_17), .E(n6402), .C(wclk), .QN(n703) );
  DFE1 \mem_reg_226][16  ( .D(D_16), .E(n6402), .C(wclk), .QN(n704) );
  DFE1 \mem_reg_226][15  ( .D(D_15), .E(n6402), .C(wclk), .QN(n705) );
  DFE1 \mem_reg_226][14  ( .D(D_14), .E(n6402), .C(wclk), .QN(n706) );
  DFE1 \mem_reg_226][13  ( .D(D_13), .E(n6402), .C(wclk), .QN(n707) );
  DFE1 \mem_reg_226][12  ( .D(D_12), .E(n6402), .C(wclk), .QN(n708) );
  DFE1 \mem_reg_226][11  ( .D(D_11), .E(n6402), .C(wclk), .QN(n709) );
  DFE1 \mem_reg_226][10  ( .D(D_10), .E(n6402), .C(wclk), .QN(n710) );
  DFE1 \mem_reg_226][9  ( .D(D_9), .E(n6402), .C(wclk), .QN(n711) );
  DFE1 \mem_reg_226][8  ( .D(D_8), .E(n6402), .C(wclk), .QN(n712) );
  DFE1 \mem_reg_226][7  ( .D(D_7), .E(n6402), .C(wclk), .QN(n713) );
  DFE1 \mem_reg_226][6  ( .D(D_6), .E(n6402), .C(wclk), .QN(n714) );
  DFE1 \mem_reg_226][5  ( .D(D_5), .E(n6402), .C(wclk), .QN(n715) );
  DFE1 \mem_reg_226][4  ( .D(D_4), .E(n6402), .C(wclk), .QN(n716) );
  DFE1 \mem_reg_226][3  ( .D(D_3), .E(n6402), .C(wclk), .QN(n717) );
  DFE1 \mem_reg_226][2  ( .D(D_2), .E(n6402), .C(wclk), .QN(n718) );
  DFE1 \mem_reg_226][1  ( .D(D_1), .E(n6402), .C(wclk), .QN(n719) );
  DFE1 \mem_reg_226][0  ( .D(D_0), .E(n6402), .C(wclk), .QN(n720) );
  DFE1 \mem_reg_225][23  ( .D(D_23), .E(n6401), .C(wclk), .QN(n721) );
  DFE1 \mem_reg_225][22  ( .D(D_22), .E(n6401), .C(wclk), .QN(n722) );
  DFE1 \mem_reg_225][21  ( .D(D_21), .E(n6401), .C(wclk), .QN(n723) );
  DFE1 \mem_reg_225][20  ( .D(D_20), .E(n6401), .C(wclk), .QN(n724) );
  DFE1 \mem_reg_225][19  ( .D(D_19), .E(n6401), .C(wclk), .QN(n725) );
  DFE1 \mem_reg_225][18  ( .D(D_18), .E(n6401), .C(wclk), .QN(n726) );
  DFE1 \mem_reg_225][17  ( .D(D_17), .E(n6401), .C(wclk), .QN(n727) );
  DFE1 \mem_reg_225][16  ( .D(D_16), .E(n6401), .C(wclk), .QN(n728) );
  DFE1 \mem_reg_225][15  ( .D(D_15), .E(n6401), .C(wclk), .QN(n729) );
  DFE1 \mem_reg_225][14  ( .D(D_14), .E(n6401), .C(wclk), .QN(n730) );
  DFE1 \mem_reg_225][13  ( .D(D_13), .E(n6401), .C(wclk), .QN(n731) );
  DFE1 \mem_reg_225][12  ( .D(D_12), .E(n6401), .C(wclk), .QN(n732) );
  DFE1 \mem_reg_225][11  ( .D(D_11), .E(n6401), .C(wclk), .QN(n733) );
  DFE1 \mem_reg_225][10  ( .D(D_10), .E(n6401), .C(wclk), .QN(n734) );
  DFE1 \mem_reg_225][9  ( .D(D_9), .E(n6401), .C(wclk), .QN(n735) );
  DFE1 \mem_reg_225][8  ( .D(D_8), .E(n6401), .C(wclk), .QN(n736) );
  DFE1 \mem_reg_225][7  ( .D(D_7), .E(n6401), .C(wclk), .QN(n737) );
  DFE1 \mem_reg_225][6  ( .D(D_6), .E(n6401), .C(wclk), .QN(n738) );
  DFE1 \mem_reg_225][5  ( .D(D_5), .E(n6401), .C(wclk), .QN(n739) );
  DFE1 \mem_reg_225][4  ( .D(D_4), .E(n6401), .C(wclk), .QN(n740) );
  DFE1 \mem_reg_225][3  ( .D(D_3), .E(n6401), .C(wclk), .QN(n741) );
  DFE1 \mem_reg_225][2  ( .D(D_2), .E(n6401), .C(wclk), .QN(n742) );
  DFE1 \mem_reg_225][1  ( .D(D_1), .E(n6401), .C(wclk), .QN(n743) );
  DFE1 \mem_reg_225][0  ( .D(D_0), .E(n6401), .C(wclk), .QN(n744) );
  DFE1 \mem_reg_224][23  ( .D(D_23), .E(n6399), .C(wclk), .QN(n745) );
  DFE1 \mem_reg_224][22  ( .D(D_22), .E(n6399), .C(wclk), .QN(n746) );
  DFE1 \mem_reg_224][21  ( .D(D_21), .E(n6399), .C(wclk), .QN(n747) );
  DFE1 \mem_reg_224][20  ( .D(D_20), .E(n6399), .C(wclk), .QN(n748) );
  DFE1 \mem_reg_224][19  ( .D(D_19), .E(n6399), .C(wclk), .QN(n749) );
  DFE1 \mem_reg_224][18  ( .D(D_18), .E(n6399), .C(wclk), .QN(n750) );
  DFE1 \mem_reg_224][17  ( .D(D_17), .E(n6399), .C(wclk), .QN(n751) );
  DFE1 \mem_reg_224][16  ( .D(D_16), .E(n6399), .C(wclk), .QN(n752) );
  DFE1 \mem_reg_224][15  ( .D(D_15), .E(n6399), .C(wclk), .QN(n753) );
  DFE1 \mem_reg_224][14  ( .D(D_14), .E(n6399), .C(wclk), .QN(n754) );
  DFE1 \mem_reg_224][13  ( .D(D_13), .E(n6399), .C(wclk), .QN(n755) );
  DFE1 \mem_reg_224][12  ( .D(D_12), .E(n6399), .C(wclk), .QN(n756) );
  DFE1 \mem_reg_224][11  ( .D(D_11), .E(n6399), .C(wclk), .QN(n757) );
  DFE1 \mem_reg_224][10  ( .D(D_10), .E(n6399), .C(wclk), .QN(n758) );
  DFE1 \mem_reg_224][9  ( .D(D_9), .E(n6399), .C(wclk), .QN(n759) );
  DFE1 \mem_reg_224][8  ( .D(D_8), .E(n6399), .C(wclk), .QN(n760) );
  DFE1 \mem_reg_224][7  ( .D(D_7), .E(n6399), .C(wclk), .QN(n761) );
  DFE1 \mem_reg_224][6  ( .D(D_6), .E(n6399), .C(wclk), .QN(n762) );
  DFE1 \mem_reg_224][5  ( .D(D_5), .E(n6399), .C(wclk), .QN(n763) );
  DFE1 \mem_reg_224][4  ( .D(D_4), .E(n6399), .C(wclk), .QN(n764) );
  DFE1 \mem_reg_224][3  ( .D(D_3), .E(n6399), .C(wclk), .QN(n765) );
  DFE1 \mem_reg_224][2  ( .D(D_2), .E(n6399), .C(wclk), .QN(n766) );
  DFE1 \mem_reg_224][1  ( .D(D_1), .E(n6399), .C(wclk), .QN(n767) );
  DFE1 \mem_reg_224][0  ( .D(D_0), .E(n6399), .C(wclk), .QN(n768) );
  DFE1 \mem_reg_223][23  ( .D(D_23), .E(n6398), .C(wclk), .QN(n769) );
  DFE1 \mem_reg_223][22  ( .D(D_22), .E(n6398), .C(wclk), .QN(n770) );
  DFE1 \mem_reg_223][21  ( .D(D_21), .E(n6398), .C(wclk), .QN(n771) );
  DFE1 \mem_reg_223][20  ( .D(D_20), .E(n6398), .C(wclk), .QN(n772) );
  DFE1 \mem_reg_223][19  ( .D(D_19), .E(n6398), .C(wclk), .QN(n773) );
  DFE1 \mem_reg_223][18  ( .D(D_18), .E(n6398), .C(wclk), .QN(n774) );
  DFE1 \mem_reg_223][17  ( .D(D_17), .E(n6398), .C(wclk), .QN(n775) );
  DFE1 \mem_reg_223][16  ( .D(D_16), .E(n6398), .C(wclk), .QN(n776) );
  DFE1 \mem_reg_223][15  ( .D(D_15), .E(n6398), .C(wclk), .QN(n777) );
  DFE1 \mem_reg_223][14  ( .D(D_14), .E(n6398), .C(wclk), .QN(n778) );
  DFE1 \mem_reg_223][13  ( .D(D_13), .E(n6398), .C(wclk), .QN(n779) );
  DFE1 \mem_reg_223][12  ( .D(D_12), .E(n6398), .C(wclk), .QN(n780) );
  DFE1 \mem_reg_223][11  ( .D(D_11), .E(n6398), .C(wclk), .QN(n781) );
  DFE1 \mem_reg_223][10  ( .D(D_10), .E(n6398), .C(wclk), .QN(n782) );
  DFE1 \mem_reg_223][9  ( .D(D_9), .E(n6398), .C(wclk), .QN(n783) );
  DFE1 \mem_reg_223][8  ( .D(D_8), .E(n6398), .C(wclk), .QN(n784) );
  DFE1 \mem_reg_223][7  ( .D(D_7), .E(n6398), .C(wclk), .QN(n785) );
  DFE1 \mem_reg_223][6  ( .D(D_6), .E(n6398), .C(wclk), .QN(n786) );
  DFE1 \mem_reg_223][5  ( .D(D_5), .E(n6398), .C(wclk), .QN(n787) );
  DFE1 \mem_reg_223][4  ( .D(D_4), .E(n6398), .C(wclk), .QN(n788) );
  DFE1 \mem_reg_223][3  ( .D(D_3), .E(n6398), .C(wclk), .QN(n789) );
  DFE1 \mem_reg_223][2  ( .D(D_2), .E(n6398), .C(wclk), .QN(n790) );
  DFE1 \mem_reg_223][1  ( .D(D_1), .E(n6398), .C(wclk), .QN(n791) );
  DFE1 \mem_reg_223][0  ( .D(D_0), .E(n6398), .C(wclk), .QN(n792) );
  DFE1 \mem_reg_222][23  ( .D(D_23), .E(n6397), .C(wclk), .QN(n793) );
  DFE1 \mem_reg_222][22  ( .D(D_22), .E(n6397), .C(wclk), .QN(n794) );
  DFE1 \mem_reg_222][21  ( .D(D_21), .E(n6397), .C(wclk), .QN(n795) );
  DFE1 \mem_reg_222][20  ( .D(D_20), .E(n6397), .C(wclk), .QN(n796) );
  DFE1 \mem_reg_222][19  ( .D(D_19), .E(n6397), .C(wclk), .QN(n797) );
  DFE1 \mem_reg_222][18  ( .D(D_18), .E(n6397), .C(wclk), .QN(n798) );
  DFE1 \mem_reg_222][17  ( .D(D_17), .E(n6397), .C(wclk), .QN(n799) );
  DFE1 \mem_reg_222][16  ( .D(D_16), .E(n6397), .C(wclk), .QN(n800) );
  DFE1 \mem_reg_222][15  ( .D(D_15), .E(n6397), .C(wclk), .QN(n801) );
  DFE1 \mem_reg_222][14  ( .D(D_14), .E(n6397), .C(wclk), .QN(n802) );
  DFE1 \mem_reg_222][13  ( .D(D_13), .E(n6397), .C(wclk), .QN(n803) );
  DFE1 \mem_reg_222][12  ( .D(D_12), .E(n6397), .C(wclk), .QN(n804) );
  DFE1 \mem_reg_222][11  ( .D(D_11), .E(n6397), .C(wclk), .QN(n805) );
  DFE1 \mem_reg_222][10  ( .D(D_10), .E(n6397), .C(wclk), .QN(n806) );
  DFE1 \mem_reg_222][9  ( .D(D_9), .E(n6397), .C(wclk), .QN(n807) );
  DFE1 \mem_reg_222][8  ( .D(D_8), .E(n6397), .C(wclk), .QN(n808) );
  DFE1 \mem_reg_222][7  ( .D(D_7), .E(n6397), .C(wclk), .QN(n809) );
  DFE1 \mem_reg_222][6  ( .D(D_6), .E(n6397), .C(wclk), .QN(n810) );
  DFE1 \mem_reg_222][5  ( .D(D_5), .E(n6397), .C(wclk), .QN(n811) );
  DFE1 \mem_reg_222][4  ( .D(D_4), .E(n6397), .C(wclk), .QN(n812) );
  DFE1 \mem_reg_222][3  ( .D(D_3), .E(n6397), .C(wclk), .QN(n813) );
  DFE1 \mem_reg_222][2  ( .D(D_2), .E(n6397), .C(wclk), .QN(n814) );
  DFE1 \mem_reg_222][1  ( .D(D_1), .E(n6397), .C(wclk), .QN(n815) );
  DFE1 \mem_reg_222][0  ( .D(D_0), .E(n6397), .C(wclk), .QN(n816) );
  DFE1 \mem_reg_221][23  ( .D(D_23), .E(n6396), .C(wclk), .QN(n817) );
  DFE1 \mem_reg_221][22  ( .D(D_22), .E(n6396), .C(wclk), .QN(n818) );
  DFE1 \mem_reg_221][21  ( .D(D_21), .E(n6396), .C(wclk), .QN(n819) );
  DFE1 \mem_reg_221][20  ( .D(D_20), .E(n6396), .C(wclk), .QN(n820) );
  DFE1 \mem_reg_221][19  ( .D(D_19), .E(n6396), .C(wclk), .QN(n821) );
  DFE1 \mem_reg_221][18  ( .D(D_18), .E(n6396), .C(wclk), .QN(n822) );
  DFE1 \mem_reg_221][17  ( .D(D_17), .E(n6396), .C(wclk), .QN(n823) );
  DFE1 \mem_reg_221][16  ( .D(D_16), .E(n6396), .C(wclk), .QN(n824) );
  DFE1 \mem_reg_221][15  ( .D(D_15), .E(n6396), .C(wclk), .QN(n825) );
  DFE1 \mem_reg_221][14  ( .D(D_14), .E(n6396), .C(wclk), .QN(n826) );
  DFE1 \mem_reg_221][13  ( .D(D_13), .E(n6396), .C(wclk), .QN(n827) );
  DFE1 \mem_reg_221][12  ( .D(D_12), .E(n6396), .C(wclk), .QN(n828) );
  DFE1 \mem_reg_221][11  ( .D(D_11), .E(n6396), .C(wclk), .QN(n829) );
  DFE1 \mem_reg_221][10  ( .D(D_10), .E(n6396), .C(wclk), .QN(n830) );
  DFE1 \mem_reg_221][9  ( .D(D_9), .E(n6396), .C(wclk), .QN(n831) );
  DFE1 \mem_reg_221][8  ( .D(D_8), .E(n6396), .C(wclk), .QN(n832) );
  DFE1 \mem_reg_221][7  ( .D(D_7), .E(n6396), .C(wclk), .QN(n833) );
  DFE1 \mem_reg_221][6  ( .D(D_6), .E(n6396), .C(wclk), .QN(n834) );
  DFE1 \mem_reg_221][5  ( .D(D_5), .E(n6396), .C(wclk), .QN(n835) );
  DFE1 \mem_reg_221][4  ( .D(D_4), .E(n6396), .C(wclk), .QN(n836) );
  DFE1 \mem_reg_221][3  ( .D(D_3), .E(n6396), .C(wclk), .QN(n837) );
  DFE1 \mem_reg_221][2  ( .D(D_2), .E(n6396), .C(wclk), .QN(n838) );
  DFE1 \mem_reg_221][1  ( .D(D_1), .E(n6396), .C(wclk), .QN(n839) );
  DFE1 \mem_reg_221][0  ( .D(D_0), .E(n6396), .C(wclk), .QN(n840) );
  DFE1 \mem_reg_220][23  ( .D(D_23), .E(n6395), .C(wclk), .QN(n841) );
  DFE1 \mem_reg_220][22  ( .D(D_22), .E(n6395), .C(wclk), .QN(n842) );
  DFE1 \mem_reg_220][21  ( .D(D_21), .E(n6395), .C(wclk), .QN(n843) );
  DFE1 \mem_reg_220][20  ( .D(D_20), .E(n6395), .C(wclk), .QN(n844) );
  DFE1 \mem_reg_220][19  ( .D(D_19), .E(n6395), .C(wclk), .QN(n845) );
  DFE1 \mem_reg_220][18  ( .D(D_18), .E(n6395), .C(wclk), .QN(n846) );
  DFE1 \mem_reg_220][17  ( .D(D_17), .E(n6395), .C(wclk), .QN(n847) );
  DFE1 \mem_reg_220][16  ( .D(D_16), .E(n6395), .C(wclk), .QN(n848) );
  DFE1 \mem_reg_220][15  ( .D(D_15), .E(n6395), .C(wclk), .QN(n849) );
  DFE1 \mem_reg_220][14  ( .D(D_14), .E(n6395), .C(wclk), .QN(n850) );
  DFE1 \mem_reg_220][13  ( .D(D_13), .E(n6395), .C(wclk), .QN(n851) );
  DFE1 \mem_reg_220][12  ( .D(D_12), .E(n6395), .C(wclk), .QN(n852) );
  DFE1 \mem_reg_220][11  ( .D(D_11), .E(n6395), .C(wclk), .QN(n853) );
  DFE1 \mem_reg_220][10  ( .D(D_10), .E(n6395), .C(wclk), .QN(n854) );
  DFE1 \mem_reg_220][9  ( .D(D_9), .E(n6395), .C(wclk), .QN(n855) );
  DFE1 \mem_reg_220][8  ( .D(D_8), .E(n6395), .C(wclk), .QN(n856) );
  DFE1 \mem_reg_220][7  ( .D(D_7), .E(n6395), .C(wclk), .QN(n857) );
  DFE1 \mem_reg_220][6  ( .D(D_6), .E(n6395), .C(wclk), .QN(n858) );
  DFE1 \mem_reg_220][5  ( .D(D_5), .E(n6395), .C(wclk), .QN(n859) );
  DFE1 \mem_reg_220][4  ( .D(D_4), .E(n6395), .C(wclk), .QN(n860) );
  DFE1 \mem_reg_220][3  ( .D(D_3), .E(n6395), .C(wclk), .QN(n861) );
  DFE1 \mem_reg_220][2  ( .D(D_2), .E(n6395), .C(wclk), .QN(n862) );
  DFE1 \mem_reg_220][1  ( .D(D_1), .E(n6395), .C(wclk), .QN(n863) );
  DFE1 \mem_reg_220][0  ( .D(D_0), .E(n6395), .C(wclk), .QN(n864) );
  DFE1 \mem_reg_219][23  ( .D(D_23), .E(n6394), .C(wclk), .QN(n865) );
  DFE1 \mem_reg_219][22  ( .D(D_22), .E(n6394), .C(wclk), .QN(n866) );
  DFE1 \mem_reg_219][21  ( .D(D_21), .E(n6394), .C(wclk), .QN(n867) );
  DFE1 \mem_reg_219][20  ( .D(D_20), .E(n6394), .C(wclk), .QN(n868) );
  DFE1 \mem_reg_219][19  ( .D(D_19), .E(n6394), .C(wclk), .QN(n869) );
  DFE1 \mem_reg_219][18  ( .D(D_18), .E(n6394), .C(wclk), .QN(n870) );
  DFE1 \mem_reg_219][17  ( .D(D_17), .E(n6394), .C(wclk), .QN(n871) );
  DFE1 \mem_reg_219][16  ( .D(D_16), .E(n6394), .C(wclk), .QN(n872) );
  DFE1 \mem_reg_219][15  ( .D(D_15), .E(n6394), .C(wclk), .QN(n873) );
  DFE1 \mem_reg_219][14  ( .D(D_14), .E(n6394), .C(wclk), .QN(n874) );
  DFE1 \mem_reg_219][13  ( .D(D_13), .E(n6394), .C(wclk), .QN(n875) );
  DFE1 \mem_reg_219][12  ( .D(D_12), .E(n6394), .C(wclk), .QN(n876) );
  DFE1 \mem_reg_219][11  ( .D(D_11), .E(n6394), .C(wclk), .QN(n877) );
  DFE1 \mem_reg_219][10  ( .D(D_10), .E(n6394), .C(wclk), .QN(n878) );
  DFE1 \mem_reg_219][9  ( .D(D_9), .E(n6394), .C(wclk), .QN(n879) );
  DFE1 \mem_reg_219][8  ( .D(D_8), .E(n6394), .C(wclk), .QN(n880) );
  DFE1 \mem_reg_219][7  ( .D(D_7), .E(n6394), .C(wclk), .QN(n881) );
  DFE1 \mem_reg_219][6  ( .D(D_6), .E(n6394), .C(wclk), .QN(n882) );
  DFE1 \mem_reg_219][5  ( .D(D_5), .E(n6394), .C(wclk), .QN(n883) );
  DFE1 \mem_reg_219][4  ( .D(D_4), .E(n6394), .C(wclk), .QN(n884) );
  DFE1 \mem_reg_219][3  ( .D(D_3), .E(n6394), .C(wclk), .QN(n885) );
  DFE1 \mem_reg_219][2  ( .D(D_2), .E(n6394), .C(wclk), .QN(n886) );
  DFE1 \mem_reg_219][1  ( .D(D_1), .E(n6394), .C(wclk), .QN(n887) );
  DFE1 \mem_reg_219][0  ( .D(D_0), .E(n6394), .C(wclk), .QN(n888) );
  DFE1 \mem_reg_218][23  ( .D(D_23), .E(n6393), .C(wclk), .QN(n889) );
  DFE1 \mem_reg_218][22  ( .D(D_22), .E(n6393), .C(wclk), .QN(n890) );
  DFE1 \mem_reg_218][21  ( .D(D_21), .E(n6393), .C(wclk), .QN(n891) );
  DFE1 \mem_reg_218][20  ( .D(D_20), .E(n6393), .C(wclk), .QN(n892) );
  DFE1 \mem_reg_218][19  ( .D(D_19), .E(n6393), .C(wclk), .QN(n893) );
  DFE1 \mem_reg_218][18  ( .D(D_18), .E(n6393), .C(wclk), .QN(n894) );
  DFE1 \mem_reg_218][17  ( .D(D_17), .E(n6393), .C(wclk), .QN(n895) );
  DFE1 \mem_reg_218][16  ( .D(D_16), .E(n6393), .C(wclk), .QN(n896) );
  DFE1 \mem_reg_218][15  ( .D(D_15), .E(n6393), .C(wclk), .QN(n897) );
  DFE1 \mem_reg_218][14  ( .D(D_14), .E(n6393), .C(wclk), .QN(n898) );
  DFE1 \mem_reg_218][13  ( .D(D_13), .E(n6393), .C(wclk), .QN(n899) );
  DFE1 \mem_reg_218][12  ( .D(D_12), .E(n6393), .C(wclk), .QN(n900) );
  DFE1 \mem_reg_218][11  ( .D(D_11), .E(n6393), .C(wclk), .QN(n901) );
  DFE1 \mem_reg_218][10  ( .D(D_10), .E(n6393), .C(wclk), .QN(n902) );
  DFE1 \mem_reg_218][9  ( .D(D_9), .E(n6393), .C(wclk), .QN(n903) );
  DFE1 \mem_reg_218][8  ( .D(D_8), .E(n6393), .C(wclk), .QN(n904) );
  DFE1 \mem_reg_218][7  ( .D(D_7), .E(n6393), .C(wclk), .QN(n905) );
  DFE1 \mem_reg_218][6  ( .D(D_6), .E(n6393), .C(wclk), .QN(n906) );
  DFE1 \mem_reg_218][5  ( .D(D_5), .E(n6393), .C(wclk), .QN(n907) );
  DFE1 \mem_reg_218][4  ( .D(D_4), .E(n6393), .C(wclk), .QN(n908) );
  DFE1 \mem_reg_218][3  ( .D(D_3), .E(n6393), .C(wclk), .QN(n909) );
  DFE1 \mem_reg_218][2  ( .D(D_2), .E(n6393), .C(wclk), .QN(n910) );
  DFE1 \mem_reg_218][1  ( .D(D_1), .E(n6393), .C(wclk), .QN(n911) );
  DFE1 \mem_reg_218][0  ( .D(D_0), .E(n6393), .C(wclk), .QN(n912) );
  DFE1 \mem_reg_217][23  ( .D(D_23), .E(n6392), .C(wclk), .QN(n913) );
  DFE1 \mem_reg_217][22  ( .D(D_22), .E(n6392), .C(wclk), .QN(n914) );
  DFE1 \mem_reg_217][21  ( .D(D_21), .E(n6392), .C(wclk), .QN(n915) );
  DFE1 \mem_reg_217][20  ( .D(D_20), .E(n6392), .C(wclk), .QN(n916) );
  DFE1 \mem_reg_217][19  ( .D(D_19), .E(n6392), .C(wclk), .QN(n917) );
  DFE1 \mem_reg_217][18  ( .D(D_18), .E(n6392), .C(wclk), .QN(n918) );
  DFE1 \mem_reg_217][17  ( .D(D_17), .E(n6392), .C(wclk), .QN(n919) );
  DFE1 \mem_reg_217][16  ( .D(D_16), .E(n6392), .C(wclk), .QN(n920) );
  DFE1 \mem_reg_217][15  ( .D(D_15), .E(n6392), .C(wclk), .QN(n921) );
  DFE1 \mem_reg_217][14  ( .D(D_14), .E(n6392), .C(wclk), .QN(n922) );
  DFE1 \mem_reg_217][13  ( .D(D_13), .E(n6392), .C(wclk), .QN(n923) );
  DFE1 \mem_reg_217][12  ( .D(D_12), .E(n6392), .C(wclk), .QN(n924) );
  DFE1 \mem_reg_217][11  ( .D(D_11), .E(n6392), .C(wclk), .QN(n925) );
  DFE1 \mem_reg_217][10  ( .D(D_10), .E(n6392), .C(wclk), .QN(n926) );
  DFE1 \mem_reg_217][9  ( .D(D_9), .E(n6392), .C(wclk), .QN(n927) );
  DFE1 \mem_reg_217][8  ( .D(D_8), .E(n6392), .C(wclk), .QN(n928) );
  DFE1 \mem_reg_217][7  ( .D(D_7), .E(n6392), .C(wclk), .QN(n929) );
  DFE1 \mem_reg_217][6  ( .D(D_6), .E(n6392), .C(wclk), .QN(n930) );
  DFE1 \mem_reg_217][5  ( .D(D_5), .E(n6392), .C(wclk), .QN(n931) );
  DFE1 \mem_reg_217][4  ( .D(D_4), .E(n6392), .C(wclk), .QN(n932) );
  DFE1 \mem_reg_217][3  ( .D(D_3), .E(n6392), .C(wclk), .QN(n933) );
  DFE1 \mem_reg_217][2  ( .D(D_2), .E(n6392), .C(wclk), .QN(n934) );
  DFE1 \mem_reg_217][1  ( .D(D_1), .E(n6392), .C(wclk), .QN(n935) );
  DFE1 \mem_reg_217][0  ( .D(D_0), .E(n6392), .C(wclk), .QN(n936) );
  DFE1 \mem_reg_216][23  ( .D(D_23), .E(n6391), .C(wclk), .QN(n937) );
  DFE1 \mem_reg_216][22  ( .D(D_22), .E(n6391), .C(wclk), .QN(n938) );
  DFE1 \mem_reg_216][21  ( .D(D_21), .E(n6391), .C(wclk), .QN(n939) );
  DFE1 \mem_reg_216][20  ( .D(D_20), .E(n6391), .C(wclk), .QN(n940) );
  DFE1 \mem_reg_216][19  ( .D(D_19), .E(n6391), .C(wclk), .QN(n941) );
  DFE1 \mem_reg_216][18  ( .D(D_18), .E(n6391), .C(wclk), .QN(n942) );
  DFE1 \mem_reg_216][17  ( .D(D_17), .E(n6391), .C(wclk), .QN(n943) );
  DFE1 \mem_reg_216][16  ( .D(D_16), .E(n6391), .C(wclk), .QN(n944) );
  DFE1 \mem_reg_216][15  ( .D(D_15), .E(n6391), .C(wclk), .QN(n945) );
  DFE1 \mem_reg_216][14  ( .D(D_14), .E(n6391), .C(wclk), .QN(n946) );
  DFE1 \mem_reg_216][13  ( .D(D_13), .E(n6391), .C(wclk), .QN(n947) );
  DFE1 \mem_reg_216][12  ( .D(D_12), .E(n6391), .C(wclk), .QN(n948) );
  DFE1 \mem_reg_216][11  ( .D(D_11), .E(n6391), .C(wclk), .QN(n949) );
  DFE1 \mem_reg_216][10  ( .D(D_10), .E(n6391), .C(wclk), .QN(n950) );
  DFE1 \mem_reg_216][9  ( .D(D_9), .E(n6391), .C(wclk), .QN(n951) );
  DFE1 \mem_reg_216][8  ( .D(D_8), .E(n6391), .C(wclk), .QN(n952) );
  DFE1 \mem_reg_216][7  ( .D(D_7), .E(n6391), .C(wclk), .QN(n953) );
  DFE1 \mem_reg_216][6  ( .D(D_6), .E(n6391), .C(wclk), .QN(n954) );
  DFE1 \mem_reg_216][5  ( .D(D_5), .E(n6391), .C(wclk), .QN(n955) );
  DFE1 \mem_reg_216][4  ( .D(D_4), .E(n6391), .C(wclk), .QN(n956) );
  DFE1 \mem_reg_216][3  ( .D(D_3), .E(n6391), .C(wclk), .QN(n957) );
  DFE1 \mem_reg_216][2  ( .D(D_2), .E(n6391), .C(wclk), .QN(n958) );
  DFE1 \mem_reg_216][1  ( .D(D_1), .E(n6391), .C(wclk), .QN(n959) );
  DFE1 \mem_reg_216][0  ( .D(D_0), .E(n6391), .C(wclk), .QN(n960) );
  DFE1 \mem_reg_215][23  ( .D(D_23), .E(n6390), .C(wclk), .QN(n961) );
  DFE1 \mem_reg_215][22  ( .D(D_22), .E(n6390), .C(wclk), .QN(n962) );
  DFE1 \mem_reg_215][21  ( .D(D_21), .E(n6390), .C(wclk), .QN(n963) );
  DFE1 \mem_reg_215][20  ( .D(D_20), .E(n6390), .C(wclk), .QN(n964) );
  DFE1 \mem_reg_215][19  ( .D(D_19), .E(n6390), .C(wclk), .QN(n965) );
  DFE1 \mem_reg_215][18  ( .D(D_18), .E(n6390), .C(wclk), .QN(n966) );
  DFE1 \mem_reg_215][17  ( .D(D_17), .E(n6390), .C(wclk), .QN(n967) );
  DFE1 \mem_reg_215][16  ( .D(D_16), .E(n6390), .C(wclk), .QN(n968) );
  DFE1 \mem_reg_215][15  ( .D(D_15), .E(n6390), .C(wclk), .QN(n969) );
  DFE1 \mem_reg_215][14  ( .D(D_14), .E(n6390), .C(wclk), .QN(n970) );
  DFE1 \mem_reg_215][13  ( .D(D_13), .E(n6390), .C(wclk), .QN(n971) );
  DFE1 \mem_reg_215][12  ( .D(D_12), .E(n6390), .C(wclk), .QN(n972) );
  DFE1 \mem_reg_215][11  ( .D(D_11), .E(n6390), .C(wclk), .QN(n973) );
  DFE1 \mem_reg_215][10  ( .D(D_10), .E(n6390), .C(wclk), .QN(n974) );
  DFE1 \mem_reg_215][9  ( .D(D_9), .E(n6390), .C(wclk), .QN(n975) );
  DFE1 \mem_reg_215][8  ( .D(D_8), .E(n6390), .C(wclk), .QN(n976) );
  DFE1 \mem_reg_215][7  ( .D(D_7), .E(n6390), .C(wclk), .QN(n977) );
  DFE1 \mem_reg_215][6  ( .D(D_6), .E(n6390), .C(wclk), .QN(n978) );
  DFE1 \mem_reg_215][5  ( .D(D_5), .E(n6390), .C(wclk), .QN(n979) );
  DFE1 \mem_reg_215][4  ( .D(D_4), .E(n6390), .C(wclk), .QN(n980) );
  DFE1 \mem_reg_215][3  ( .D(D_3), .E(n6390), .C(wclk), .QN(n981) );
  DFE1 \mem_reg_215][2  ( .D(D_2), .E(n6390), .C(wclk), .QN(n982) );
  DFE1 \mem_reg_215][1  ( .D(D_1), .E(n6390), .C(wclk), .QN(n983) );
  DFE1 \mem_reg_215][0  ( .D(D_0), .E(n6390), .C(wclk), .QN(n984) );
  DFE1 \mem_reg_214][23  ( .D(D_23), .E(n6389), .C(wclk), .QN(n985) );
  DFE1 \mem_reg_214][22  ( .D(D_22), .E(n6389), .C(wclk), .QN(n986) );
  DFE1 \mem_reg_214][21  ( .D(D_21), .E(n6389), .C(wclk), .QN(n987) );
  DFE1 \mem_reg_214][20  ( .D(D_20), .E(n6389), .C(wclk), .QN(n988) );
  DFE1 \mem_reg_214][19  ( .D(D_19), .E(n6389), .C(wclk), .QN(n989) );
  DFE1 \mem_reg_214][18  ( .D(D_18), .E(n6389), .C(wclk), .QN(n990) );
  DFE1 \mem_reg_214][17  ( .D(D_17), .E(n6389), .C(wclk), .QN(n991) );
  DFE1 \mem_reg_214][16  ( .D(D_16), .E(n6389), .C(wclk), .QN(n992) );
  DFE1 \mem_reg_214][15  ( .D(D_15), .E(n6389), .C(wclk), .QN(n993) );
  DFE1 \mem_reg_214][14  ( .D(D_14), .E(n6389), .C(wclk), .QN(n994) );
  DFE1 \mem_reg_214][13  ( .D(D_13), .E(n6389), .C(wclk), .QN(n995) );
  DFE1 \mem_reg_214][12  ( .D(D_12), .E(n6389), .C(wclk), .QN(n996) );
  DFE1 \mem_reg_214][11  ( .D(D_11), .E(n6389), .C(wclk), .QN(n997) );
  DFE1 \mem_reg_214][10  ( .D(D_10), .E(n6389), .C(wclk), .QN(n998) );
  DFE1 \mem_reg_214][9  ( .D(D_9), .E(n6389), .C(wclk), .QN(n999) );
  DFE1 \mem_reg_214][8  ( .D(D_8), .E(n6389), .C(wclk), .QN(n1000) );
  DFE1 \mem_reg_214][7  ( .D(D_7), .E(n6389), .C(wclk), .QN(n1001) );
  DFE1 \mem_reg_214][6  ( .D(D_6), .E(n6389), .C(wclk), .QN(n1002) );
  DFE1 \mem_reg_214][5  ( .D(D_5), .E(n6389), .C(wclk), .QN(n1003) );
  DFE1 \mem_reg_214][4  ( .D(D_4), .E(n6389), .C(wclk), .QN(n1004) );
  DFE1 \mem_reg_214][3  ( .D(D_3), .E(n6389), .C(wclk), .QN(n1005) );
  DFE1 \mem_reg_214][2  ( .D(D_2), .E(n6389), .C(wclk), .QN(n1006) );
  DFE1 \mem_reg_214][1  ( .D(D_1), .E(n6389), .C(wclk), .QN(n1007) );
  DFE1 \mem_reg_214][0  ( .D(D_0), .E(n6389), .C(wclk), .QN(n1008) );
  DFE1 \mem_reg_213][23  ( .D(D_23), .E(n6388), .C(wclk), .QN(n1009) );
  DFE1 \mem_reg_213][22  ( .D(D_22), .E(n6388), .C(wclk), .QN(n1010) );
  DFE1 \mem_reg_213][21  ( .D(D_21), .E(n6388), .C(wclk), .QN(n1011) );
  DFE1 \mem_reg_213][20  ( .D(D_20), .E(n6388), .C(wclk), .QN(n1012) );
  DFE1 \mem_reg_213][19  ( .D(D_19), .E(n6388), .C(wclk), .QN(n1013) );
  DFE1 \mem_reg_213][18  ( .D(D_18), .E(n6388), .C(wclk), .QN(n1014) );
  DFE1 \mem_reg_213][17  ( .D(D_17), .E(n6388), .C(wclk), .QN(n1015) );
  DFE1 \mem_reg_213][16  ( .D(D_16), .E(n6388), .C(wclk), .QN(n1016) );
  DFE1 \mem_reg_213][15  ( .D(D_15), .E(n6388), .C(wclk), .QN(n1017) );
  DFE1 \mem_reg_213][14  ( .D(D_14), .E(n6388), .C(wclk), .QN(n1018) );
  DFE1 \mem_reg_213][13  ( .D(D_13), .E(n6388), .C(wclk), .QN(n1019) );
  DFE1 \mem_reg_213][12  ( .D(D_12), .E(n6388), .C(wclk), .QN(n1020) );
  DFE1 \mem_reg_213][11  ( .D(D_11), .E(n6388), .C(wclk), .QN(n1021) );
  DFE1 \mem_reg_213][10  ( .D(D_10), .E(n6388), .C(wclk), .QN(n1022) );
  DFE1 \mem_reg_213][9  ( .D(D_9), .E(n6388), .C(wclk), .QN(n1023) );
  DFE1 \mem_reg_213][8  ( .D(D_8), .E(n6388), .C(wclk), .QN(n1024) );
  DFE1 \mem_reg_213][7  ( .D(D_7), .E(n6388), .C(wclk), .QN(n1025) );
  DFE1 \mem_reg_213][6  ( .D(D_6), .E(n6388), .C(wclk), .QN(n1026) );
  DFE1 \mem_reg_213][5  ( .D(D_5), .E(n6388), .C(wclk), .QN(n1027) );
  DFE1 \mem_reg_213][4  ( .D(D_4), .E(n6388), .C(wclk), .QN(n1028) );
  DFE1 \mem_reg_213][3  ( .D(D_3), .E(n6388), .C(wclk), .QN(n1029) );
  DFE1 \mem_reg_213][2  ( .D(D_2), .E(n6388), .C(wclk), .QN(n1030) );
  DFE1 \mem_reg_213][1  ( .D(D_1), .E(n6388), .C(wclk), .QN(n1031) );
  DFE1 \mem_reg_213][0  ( .D(D_0), .E(n6388), .C(wclk), .QN(n1032) );
  DFE1 \mem_reg_212][23  ( .D(D_23), .E(n6387), .C(wclk), .QN(n1033) );
  DFE1 \mem_reg_212][22  ( .D(D_22), .E(n6387), .C(wclk), .QN(n1034) );
  DFE1 \mem_reg_212][21  ( .D(D_21), .E(n6387), .C(wclk), .QN(n1035) );
  DFE1 \mem_reg_212][20  ( .D(D_20), .E(n6387), .C(wclk), .QN(n1036) );
  DFE1 \mem_reg_212][19  ( .D(D_19), .E(n6387), .C(wclk), .QN(n1037) );
  DFE1 \mem_reg_212][18  ( .D(D_18), .E(n6387), .C(wclk), .QN(n1038) );
  DFE1 \mem_reg_212][17  ( .D(D_17), .E(n6387), .C(wclk), .QN(n1039) );
  DFE1 \mem_reg_212][16  ( .D(D_16), .E(n6387), .C(wclk), .QN(n1040) );
  DFE1 \mem_reg_212][15  ( .D(D_15), .E(n6387), .C(wclk), .QN(n1041) );
  DFE1 \mem_reg_212][14  ( .D(D_14), .E(n6387), .C(wclk), .QN(n1042) );
  DFE1 \mem_reg_212][13  ( .D(D_13), .E(n6387), .C(wclk), .QN(n1043) );
  DFE1 \mem_reg_212][12  ( .D(D_12), .E(n6387), .C(wclk), .QN(n1044) );
  DFE1 \mem_reg_212][11  ( .D(D_11), .E(n6387), .C(wclk), .QN(n1045) );
  DFE1 \mem_reg_212][10  ( .D(D_10), .E(n6387), .C(wclk), .QN(n1046) );
  DFE1 \mem_reg_212][9  ( .D(D_9), .E(n6387), .C(wclk), .QN(n1047) );
  DFE1 \mem_reg_212][8  ( .D(D_8), .E(n6387), .C(wclk), .QN(n1048) );
  DFE1 \mem_reg_212][7  ( .D(D_7), .E(n6387), .C(wclk), .QN(n1049) );
  DFE1 \mem_reg_212][6  ( .D(D_6), .E(n6387), .C(wclk), .QN(n1050) );
  DFE1 \mem_reg_212][5  ( .D(D_5), .E(n6387), .C(wclk), .QN(n1051) );
  DFE1 \mem_reg_212][4  ( .D(D_4), .E(n6387), .C(wclk), .QN(n1052) );
  DFE1 \mem_reg_212][3  ( .D(D_3), .E(n6387), .C(wclk), .QN(n1053) );
  DFE1 \mem_reg_212][2  ( .D(D_2), .E(n6387), .C(wclk), .QN(n1054) );
  DFE1 \mem_reg_212][1  ( .D(D_1), .E(n6387), .C(wclk), .QN(n1055) );
  DFE1 \mem_reg_212][0  ( .D(D_0), .E(n6387), .C(wclk), .QN(n1056) );
  DFE1 \mem_reg_211][23  ( .D(D_23), .E(n6386), .C(wclk), .QN(n1057) );
  DFE1 \mem_reg_211][22  ( .D(D_22), .E(n6386), .C(wclk), .QN(n1058) );
  DFE1 \mem_reg_211][21  ( .D(D_21), .E(n6386), .C(wclk), .QN(n1059) );
  DFE1 \mem_reg_211][20  ( .D(D_20), .E(n6386), .C(wclk), .QN(n1060) );
  DFE1 \mem_reg_211][19  ( .D(D_19), .E(n6386), .C(wclk), .QN(n1061) );
  DFE1 \mem_reg_211][18  ( .D(D_18), .E(n6386), .C(wclk), .QN(n1062) );
  DFE1 \mem_reg_211][17  ( .D(D_17), .E(n6386), .C(wclk), .QN(n1063) );
  DFE1 \mem_reg_211][16  ( .D(D_16), .E(n6386), .C(wclk), .QN(n1064) );
  DFE1 \mem_reg_211][15  ( .D(D_15), .E(n6386), .C(wclk), .QN(n1065) );
  DFE1 \mem_reg_211][14  ( .D(D_14), .E(n6386), .C(wclk), .QN(n1066) );
  DFE1 \mem_reg_211][13  ( .D(D_13), .E(n6386), .C(wclk), .QN(n1067) );
  DFE1 \mem_reg_211][12  ( .D(D_12), .E(n6386), .C(wclk), .QN(n1068) );
  DFE1 \mem_reg_211][11  ( .D(D_11), .E(n6386), .C(wclk), .QN(n1069) );
  DFE1 \mem_reg_211][10  ( .D(D_10), .E(n6386), .C(wclk), .QN(n1070) );
  DFE1 \mem_reg_211][9  ( .D(D_9), .E(n6386), .C(wclk), .QN(n1071) );
  DFE1 \mem_reg_211][8  ( .D(D_8), .E(n6386), .C(wclk), .QN(n1072) );
  DFE1 \mem_reg_211][7  ( .D(D_7), .E(n6386), .C(wclk), .QN(n1073) );
  DFE1 \mem_reg_211][6  ( .D(D_6), .E(n6386), .C(wclk), .QN(n1074) );
  DFE1 \mem_reg_211][5  ( .D(D_5), .E(n6386), .C(wclk), .QN(n1075) );
  DFE1 \mem_reg_211][4  ( .D(D_4), .E(n6386), .C(wclk), .QN(n1076) );
  DFE1 \mem_reg_211][3  ( .D(D_3), .E(n6386), .C(wclk), .QN(n1077) );
  DFE1 \mem_reg_211][2  ( .D(D_2), .E(n6386), .C(wclk), .QN(n1078) );
  DFE1 \mem_reg_211][1  ( .D(D_1), .E(n6386), .C(wclk), .QN(n1079) );
  DFE1 \mem_reg_211][0  ( .D(D_0), .E(n6386), .C(wclk), .QN(n1080) );
  DFE1 \mem_reg_210][23  ( .D(D_23), .E(n6385), .C(wclk), .QN(n1081) );
  DFE1 \mem_reg_210][22  ( .D(D_22), .E(n6385), .C(wclk), .QN(n1082) );
  DFE1 \mem_reg_210][21  ( .D(D_21), .E(n6385), .C(wclk), .QN(n1083) );
  DFE1 \mem_reg_210][20  ( .D(D_20), .E(n6385), .C(wclk), .QN(n1084) );
  DFE1 \mem_reg_210][19  ( .D(D_19), .E(n6385), .C(wclk), .QN(n1085) );
  DFE1 \mem_reg_210][18  ( .D(D_18), .E(n6385), .C(wclk), .QN(n1086) );
  DFE1 \mem_reg_210][17  ( .D(D_17), .E(n6385), .C(wclk), .QN(n1087) );
  DFE1 \mem_reg_210][16  ( .D(D_16), .E(n6385), .C(wclk), .QN(n1088) );
  DFE1 \mem_reg_210][15  ( .D(D_15), .E(n6385), .C(wclk), .QN(n1089) );
  DFE1 \mem_reg_210][14  ( .D(D_14), .E(n6385), .C(wclk), .QN(n1090) );
  DFE1 \mem_reg_210][13  ( .D(D_13), .E(n6385), .C(wclk), .QN(n1091) );
  DFE1 \mem_reg_210][12  ( .D(D_12), .E(n6385), .C(wclk), .QN(n1092) );
  DFE1 \mem_reg_210][11  ( .D(D_11), .E(n6385), .C(wclk), .QN(n1093) );
  DFE1 \mem_reg_210][10  ( .D(D_10), .E(n6385), .C(wclk), .QN(n1094) );
  DFE1 \mem_reg_210][9  ( .D(D_9), .E(n6385), .C(wclk), .QN(n1095) );
  DFE1 \mem_reg_210][8  ( .D(D_8), .E(n6385), .C(wclk), .QN(n1096) );
  DFE1 \mem_reg_210][7  ( .D(D_7), .E(n6385), .C(wclk), .QN(n1097) );
  DFE1 \mem_reg_210][6  ( .D(D_6), .E(n6385), .C(wclk), .QN(n1098) );
  DFE1 \mem_reg_210][5  ( .D(D_5), .E(n6385), .C(wclk), .QN(n1099) );
  DFE1 \mem_reg_210][4  ( .D(D_4), .E(n6385), .C(wclk), .QN(n1100) );
  DFE1 \mem_reg_210][3  ( .D(D_3), .E(n6385), .C(wclk), .QN(n1101) );
  DFE1 \mem_reg_210][2  ( .D(D_2), .E(n6385), .C(wclk), .QN(n1102) );
  DFE1 \mem_reg_210][1  ( .D(D_1), .E(n6385), .C(wclk), .QN(n1103) );
  DFE1 \mem_reg_210][0  ( .D(D_0), .E(n6385), .C(wclk), .QN(n1104) );
  DFE1 \mem_reg_209][23  ( .D(D_23), .E(n6384), .C(wclk), .QN(n1105) );
  DFE1 \mem_reg_209][22  ( .D(D_22), .E(n6384), .C(wclk), .QN(n1106) );
  DFE1 \mem_reg_209][21  ( .D(D_21), .E(n6384), .C(wclk), .QN(n1107) );
  DFE1 \mem_reg_209][20  ( .D(D_20), .E(n6384), .C(wclk), .QN(n1108) );
  DFE1 \mem_reg_209][19  ( .D(D_19), .E(n6384), .C(wclk), .QN(n1109) );
  DFE1 \mem_reg_209][18  ( .D(D_18), .E(n6384), .C(wclk), .QN(n1110) );
  DFE1 \mem_reg_209][17  ( .D(D_17), .E(n6384), .C(wclk), .QN(n1111) );
  DFE1 \mem_reg_209][16  ( .D(D_16), .E(n6384), .C(wclk), .QN(n1112) );
  DFE1 \mem_reg_209][15  ( .D(D_15), .E(n6384), .C(wclk), .QN(n1113) );
  DFE1 \mem_reg_209][14  ( .D(D_14), .E(n6384), .C(wclk), .QN(n1114) );
  DFE1 \mem_reg_209][13  ( .D(D_13), .E(n6384), .C(wclk), .QN(n1115) );
  DFE1 \mem_reg_209][12  ( .D(D_12), .E(n6384), .C(wclk), .QN(n1116) );
  DFE1 \mem_reg_209][11  ( .D(D_11), .E(n6384), .C(wclk), .QN(n1117) );
  DFE1 \mem_reg_209][10  ( .D(D_10), .E(n6384), .C(wclk), .QN(n1118) );
  DFE1 \mem_reg_209][9  ( .D(D_9), .E(n6384), .C(wclk), .QN(n1119) );
  DFE1 \mem_reg_209][8  ( .D(D_8), .E(n6384), .C(wclk), .QN(n1120) );
  DFE1 \mem_reg_209][7  ( .D(D_7), .E(n6384), .C(wclk), .QN(n1121) );
  DFE1 \mem_reg_209][6  ( .D(D_6), .E(n6384), .C(wclk), .QN(n1122) );
  DFE1 \mem_reg_209][5  ( .D(D_5), .E(n6384), .C(wclk), .QN(n1123) );
  DFE1 \mem_reg_209][4  ( .D(D_4), .E(n6384), .C(wclk), .QN(n1124) );
  DFE1 \mem_reg_209][3  ( .D(D_3), .E(n6384), .C(wclk), .QN(n1125) );
  DFE1 \mem_reg_209][2  ( .D(D_2), .E(n6384), .C(wclk), .QN(n1126) );
  DFE1 \mem_reg_209][1  ( .D(D_1), .E(n6384), .C(wclk), .QN(n1127) );
  DFE1 \mem_reg_209][0  ( .D(D_0), .E(n6384), .C(wclk), .QN(n1128) );
  DFE1 \mem_reg_208][23  ( .D(D_23), .E(n6382), .C(wclk), .QN(n1129) );
  DFE1 \mem_reg_208][22  ( .D(D_22), .E(n6382), .C(wclk), .QN(n1130) );
  DFE1 \mem_reg_208][21  ( .D(D_21), .E(n6382), .C(wclk), .QN(n1131) );
  DFE1 \mem_reg_208][20  ( .D(D_20), .E(n6382), .C(wclk), .QN(n1132) );
  DFE1 \mem_reg_208][19  ( .D(D_19), .E(n6382), .C(wclk), .QN(n1133) );
  DFE1 \mem_reg_208][18  ( .D(D_18), .E(n6382), .C(wclk), .QN(n1134) );
  DFE1 \mem_reg_208][17  ( .D(D_17), .E(n6382), .C(wclk), .QN(n1135) );
  DFE1 \mem_reg_208][16  ( .D(D_16), .E(n6382), .C(wclk), .QN(n1136) );
  DFE1 \mem_reg_208][15  ( .D(D_15), .E(n6382), .C(wclk), .QN(n1137) );
  DFE1 \mem_reg_208][14  ( .D(D_14), .E(n6382), .C(wclk), .QN(n1138) );
  DFE1 \mem_reg_208][13  ( .D(D_13), .E(n6382), .C(wclk), .QN(n1139) );
  DFE1 \mem_reg_208][12  ( .D(D_12), .E(n6382), .C(wclk), .QN(n1140) );
  DFE1 \mem_reg_208][11  ( .D(D_11), .E(n6382), .C(wclk), .QN(n1141) );
  DFE1 \mem_reg_208][10  ( .D(D_10), .E(n6382), .C(wclk), .QN(n1142) );
  DFE1 \mem_reg_208][9  ( .D(D_9), .E(n6382), .C(wclk), .QN(n1143) );
  DFE1 \mem_reg_208][8  ( .D(D_8), .E(n6382), .C(wclk), .QN(n1144) );
  DFE1 \mem_reg_208][7  ( .D(D_7), .E(n6382), .C(wclk), .QN(n1145) );
  DFE1 \mem_reg_208][6  ( .D(D_6), .E(n6382), .C(wclk), .QN(n1146) );
  DFE1 \mem_reg_208][5  ( .D(D_5), .E(n6382), .C(wclk), .QN(n1147) );
  DFE1 \mem_reg_208][4  ( .D(D_4), .E(n6382), .C(wclk), .QN(n1148) );
  DFE1 \mem_reg_208][3  ( .D(D_3), .E(n6382), .C(wclk), .QN(n1149) );
  DFE1 \mem_reg_208][2  ( .D(D_2), .E(n6382), .C(wclk), .QN(n1150) );
  DFE1 \mem_reg_208][1  ( .D(D_1), .E(n6382), .C(wclk), .QN(n1151) );
  DFE1 \mem_reg_208][0  ( .D(D_0), .E(n6382), .C(wclk), .QN(n1152) );
  DFE1 \mem_reg_111][23  ( .D(D_23), .E(n6273), .C(wclk), .QN(n3457) );
  DFE1 \mem_reg_111][22  ( .D(D_22), .E(n6273), .C(wclk), .QN(n3458) );
  DFE1 \mem_reg_111][21  ( .D(D_21), .E(n6273), .C(wclk), .QN(n3459) );
  DFE1 \mem_reg_111][20  ( .D(D_20), .E(n6273), .C(wclk), .QN(n3460) );
  DFE1 \mem_reg_111][19  ( .D(D_19), .E(n6273), .C(wclk), .QN(n3461) );
  DFE1 \mem_reg_111][18  ( .D(D_18), .E(n6273), .C(wclk), .QN(n3462) );
  DFE1 \mem_reg_111][17  ( .D(D_17), .E(n6273), .C(wclk), .QN(n3463) );
  DFE1 \mem_reg_111][16  ( .D(D_16), .E(n6273), .C(wclk), .QN(n3464) );
  DFE1 \mem_reg_111][15  ( .D(D_15), .E(n6273), .C(wclk), .QN(n3465) );
  DFE1 \mem_reg_111][14  ( .D(D_14), .E(n6273), .C(wclk), .QN(n3466) );
  DFE1 \mem_reg_111][13  ( .D(D_13), .E(n6273), .C(wclk), .QN(n3467) );
  DFE1 \mem_reg_111][12  ( .D(D_12), .E(n6273), .C(wclk), .QN(n3468) );
  DFE1 \mem_reg_111][11  ( .D(D_11), .E(n6273), .C(wclk), .QN(n3469) );
  DFE1 \mem_reg_111][10  ( .D(D_10), .E(n6273), .C(wclk), .QN(n3470) );
  DFE1 \mem_reg_111][9  ( .D(D_9), .E(n6273), .C(wclk), .QN(n3471) );
  DFE1 \mem_reg_111][8  ( .D(D_8), .E(n6273), .C(wclk), .QN(n3472) );
  DFE1 \mem_reg_111][7  ( .D(D_7), .E(n6273), .C(wclk), .QN(n3473) );
  DFE1 \mem_reg_111][6  ( .D(D_6), .E(n6273), .C(wclk), .QN(n3474) );
  DFE1 \mem_reg_111][5  ( .D(D_5), .E(n6273), .C(wclk), .QN(n3475) );
  DFE1 \mem_reg_111][4  ( .D(D_4), .E(n6273), .C(wclk), .QN(n3476) );
  DFE1 \mem_reg_111][3  ( .D(D_3), .E(n6273), .C(wclk), .QN(n3477) );
  DFE1 \mem_reg_111][2  ( .D(D_2), .E(n6273), .C(wclk), .QN(n3478) );
  DFE1 \mem_reg_111][1  ( .D(D_1), .E(n6273), .C(wclk), .QN(n3479) );
  DFE1 \mem_reg_111][0  ( .D(D_0), .E(n6273), .C(wclk), .QN(n3480) );
  DFE1 \mem_reg_110][23  ( .D(D_23), .E(n6272), .C(wclk), .QN(n3481) );
  DFE1 \mem_reg_110][22  ( .D(D_22), .E(n6272), .C(wclk), .QN(n3482) );
  DFE1 \mem_reg_110][21  ( .D(D_21), .E(n6272), .C(wclk), .QN(n3483) );
  DFE1 \mem_reg_110][20  ( .D(D_20), .E(n6272), .C(wclk), .QN(n3484) );
  DFE1 \mem_reg_110][19  ( .D(D_19), .E(n6272), .C(wclk), .QN(n3485) );
  DFE1 \mem_reg_110][18  ( .D(D_18), .E(n6272), .C(wclk), .QN(n3486) );
  DFE1 \mem_reg_110][17  ( .D(D_17), .E(n6272), .C(wclk), .QN(n3487) );
  DFE1 \mem_reg_110][16  ( .D(D_16), .E(n6272), .C(wclk), .QN(n3488) );
  DFE1 \mem_reg_110][15  ( .D(D_15), .E(n6272), .C(wclk), .QN(n3489) );
  DFE1 \mem_reg_110][14  ( .D(D_14), .E(n6272), .C(wclk), .QN(n3490) );
  DFE1 \mem_reg_110][13  ( .D(D_13), .E(n6272), .C(wclk), .QN(n3491) );
  DFE1 \mem_reg_110][12  ( .D(D_12), .E(n6272), .C(wclk), .QN(n3492) );
  DFE1 \mem_reg_110][11  ( .D(D_11), .E(n6272), .C(wclk), .QN(n3493) );
  DFE1 \mem_reg_110][10  ( .D(D_10), .E(n6272), .C(wclk), .QN(n3494) );
  DFE1 \mem_reg_110][9  ( .D(D_9), .E(n6272), .C(wclk), .QN(n3495) );
  DFE1 \mem_reg_110][8  ( .D(D_8), .E(n6272), .C(wclk), .QN(n3496) );
  DFE1 \mem_reg_110][7  ( .D(D_7), .E(n6272), .C(wclk), .QN(n3497) );
  DFE1 \mem_reg_110][6  ( .D(D_6), .E(n6272), .C(wclk), .QN(n3498) );
  DFE1 \mem_reg_110][5  ( .D(D_5), .E(n6272), .C(wclk), .QN(n3499) );
  DFE1 \mem_reg_110][4  ( .D(D_4), .E(n6272), .C(wclk), .QN(n3500) );
  DFE1 \mem_reg_110][3  ( .D(D_3), .E(n6272), .C(wclk), .QN(n3501) );
  DFE1 \mem_reg_110][2  ( .D(D_2), .E(n6272), .C(wclk), .QN(n3502) );
  DFE1 \mem_reg_110][1  ( .D(D_1), .E(n6272), .C(wclk), .QN(n3503) );
  DFE1 \mem_reg_110][0  ( .D(D_0), .E(n6272), .C(wclk), .QN(n3504) );
  DFE1 \mem_reg_109][23  ( .D(D_23), .E(n6271), .C(wclk), .QN(n3505) );
  DFE1 \mem_reg_109][22  ( .D(D_22), .E(n6271), .C(wclk), .QN(n3506) );
  DFE1 \mem_reg_109][21  ( .D(D_21), .E(n6271), .C(wclk), .QN(n3507) );
  DFE1 \mem_reg_109][20  ( .D(D_20), .E(n6271), .C(wclk), .QN(n3508) );
  DFE1 \mem_reg_109][19  ( .D(D_19), .E(n6271), .C(wclk), .QN(n3509) );
  DFE1 \mem_reg_109][18  ( .D(D_18), .E(n6271), .C(wclk), .QN(n3510) );
  DFE1 \mem_reg_109][17  ( .D(D_17), .E(n6271), .C(wclk), .QN(n3511) );
  DFE1 \mem_reg_109][16  ( .D(D_16), .E(n6271), .C(wclk), .QN(n3512) );
  DFE1 \mem_reg_109][15  ( .D(D_15), .E(n6271), .C(wclk), .QN(n3513) );
  DFE1 \mem_reg_109][14  ( .D(D_14), .E(n6271), .C(wclk), .QN(n3514) );
  DFE1 \mem_reg_109][13  ( .D(D_13), .E(n6271), .C(wclk), .QN(n3515) );
  DFE1 \mem_reg_109][12  ( .D(D_12), .E(n6271), .C(wclk), .QN(n3516) );
  DFE1 \mem_reg_109][11  ( .D(D_11), .E(n6271), .C(wclk), .QN(n3517) );
  DFE1 \mem_reg_109][10  ( .D(D_10), .E(n6271), .C(wclk), .QN(n3518) );
  DFE1 \mem_reg_109][9  ( .D(D_9), .E(n6271), .C(wclk), .QN(n3519) );
  DFE1 \mem_reg_109][8  ( .D(D_8), .E(n6271), .C(wclk), .QN(n3520) );
  DFE1 \mem_reg_109][7  ( .D(D_7), .E(n6271), .C(wclk), .QN(n3521) );
  DFE1 \mem_reg_109][6  ( .D(D_6), .E(n6271), .C(wclk), .QN(n3522) );
  DFE1 \mem_reg_109][5  ( .D(D_5), .E(n6271), .C(wclk), .QN(n3523) );
  DFE1 \mem_reg_109][4  ( .D(D_4), .E(n6271), .C(wclk), .QN(n3524) );
  DFE1 \mem_reg_109][3  ( .D(D_3), .E(n6271), .C(wclk), .QN(n3525) );
  DFE1 \mem_reg_109][2  ( .D(D_2), .E(n6271), .C(wclk), .QN(n3526) );
  DFE1 \mem_reg_109][1  ( .D(D_1), .E(n6271), .C(wclk), .QN(n3527) );
  DFE1 \mem_reg_109][0  ( .D(D_0), .E(n6271), .C(wclk), .QN(n3528) );
  DFE1 \mem_reg_108][23  ( .D(D_23), .E(n6270), .C(wclk), .QN(n3529) );
  DFE1 \mem_reg_108][22  ( .D(D_22), .E(n6270), .C(wclk), .QN(n3530) );
  DFE1 \mem_reg_108][21  ( .D(D_21), .E(n6270), .C(wclk), .QN(n3531) );
  DFE1 \mem_reg_108][20  ( .D(D_20), .E(n6270), .C(wclk), .QN(n3532) );
  DFE1 \mem_reg_108][19  ( .D(D_19), .E(n6270), .C(wclk), .QN(n3533) );
  DFE1 \mem_reg_108][18  ( .D(D_18), .E(n6270), .C(wclk), .QN(n3534) );
  DFE1 \mem_reg_108][17  ( .D(D_17), .E(n6270), .C(wclk), .QN(n3535) );
  DFE1 \mem_reg_108][16  ( .D(D_16), .E(n6270), .C(wclk), .QN(n3536) );
  DFE1 \mem_reg_108][15  ( .D(D_15), .E(n6270), .C(wclk), .QN(n3537) );
  DFE1 \mem_reg_108][14  ( .D(D_14), .E(n6270), .C(wclk), .QN(n3538) );
  DFE1 \mem_reg_108][13  ( .D(D_13), .E(n6270), .C(wclk), .QN(n3539) );
  DFE1 \mem_reg_108][12  ( .D(D_12), .E(n6270), .C(wclk), .QN(n3540) );
  DFE1 \mem_reg_108][11  ( .D(D_11), .E(n6270), .C(wclk), .QN(n3541) );
  DFE1 \mem_reg_108][10  ( .D(D_10), .E(n6270), .C(wclk), .QN(n3542) );
  DFE1 \mem_reg_108][9  ( .D(D_9), .E(n6270), .C(wclk), .QN(n3543) );
  DFE1 \mem_reg_108][8  ( .D(D_8), .E(n6270), .C(wclk), .QN(n3544) );
  DFE1 \mem_reg_108][7  ( .D(D_7), .E(n6270), .C(wclk), .QN(n3545) );
  DFE1 \mem_reg_108][6  ( .D(D_6), .E(n6270), .C(wclk), .QN(n3546) );
  DFE1 \mem_reg_108][5  ( .D(D_5), .E(n6270), .C(wclk), .QN(n3547) );
  DFE1 \mem_reg_108][4  ( .D(D_4), .E(n6270), .C(wclk), .QN(n3548) );
  DFE1 \mem_reg_108][3  ( .D(D_3), .E(n6270), .C(wclk), .QN(n3549) );
  DFE1 \mem_reg_108][2  ( .D(D_2), .E(n6270), .C(wclk), .QN(n3550) );
  DFE1 \mem_reg_108][1  ( .D(D_1), .E(n6270), .C(wclk), .QN(n3551) );
  DFE1 \mem_reg_108][0  ( .D(D_0), .E(n6270), .C(wclk), .QN(n3552) );
  DFE1 \mem_reg_107][23  ( .D(D_23), .E(n6269), .C(wclk), .QN(n3553) );
  DFE1 \mem_reg_107][22  ( .D(D_22), .E(n6269), .C(wclk), .QN(n3554) );
  DFE1 \mem_reg_107][21  ( .D(D_21), .E(n6269), .C(wclk), .QN(n3555) );
  DFE1 \mem_reg_107][20  ( .D(D_20), .E(n6269), .C(wclk), .QN(n3556) );
  DFE1 \mem_reg_107][19  ( .D(D_19), .E(n6269), .C(wclk), .QN(n3557) );
  DFE1 \mem_reg_107][18  ( .D(D_18), .E(n6269), .C(wclk), .QN(n3558) );
  DFE1 \mem_reg_107][17  ( .D(D_17), .E(n6269), .C(wclk), .QN(n3559) );
  DFE1 \mem_reg_107][16  ( .D(D_16), .E(n6269), .C(wclk), .QN(n3560) );
  DFE1 \mem_reg_107][15  ( .D(D_15), .E(n6269), .C(wclk), .QN(n3561) );
  DFE1 \mem_reg_107][14  ( .D(D_14), .E(n6269), .C(wclk), .QN(n3562) );
  DFE1 \mem_reg_107][13  ( .D(D_13), .E(n6269), .C(wclk), .QN(n3563) );
  DFE1 \mem_reg_107][12  ( .D(D_12), .E(n6269), .C(wclk), .QN(n3564) );
  DFE1 \mem_reg_107][11  ( .D(D_11), .E(n6269), .C(wclk), .QN(n3565) );
  DFE1 \mem_reg_107][10  ( .D(D_10), .E(n6269), .C(wclk), .QN(n3566) );
  DFE1 \mem_reg_107][9  ( .D(D_9), .E(n6269), .C(wclk), .QN(n3567) );
  DFE1 \mem_reg_107][8  ( .D(D_8), .E(n6269), .C(wclk), .QN(n3568) );
  DFE1 \mem_reg_107][7  ( .D(D_7), .E(n6269), .C(wclk), .QN(n3569) );
  DFE1 \mem_reg_107][6  ( .D(D_6), .E(n6269), .C(wclk), .QN(n3570) );
  DFE1 \mem_reg_107][5  ( .D(D_5), .E(n6269), .C(wclk), .QN(n3571) );
  DFE1 \mem_reg_107][4  ( .D(D_4), .E(n6269), .C(wclk), .QN(n3572) );
  DFE1 \mem_reg_107][3  ( .D(D_3), .E(n6269), .C(wclk), .QN(n3573) );
  DFE1 \mem_reg_107][2  ( .D(D_2), .E(n6269), .C(wclk), .QN(n3574) );
  DFE1 \mem_reg_107][1  ( .D(D_1), .E(n6269), .C(wclk), .QN(n3575) );
  DFE1 \mem_reg_107][0  ( .D(D_0), .E(n6269), .C(wclk), .QN(n3576) );
  DFE1 \mem_reg_106][23  ( .D(D_23), .E(n6268), .C(wclk), .QN(n3577) );
  DFE1 \mem_reg_106][22  ( .D(D_22), .E(n6268), .C(wclk), .QN(n3578) );
  DFE1 \mem_reg_106][21  ( .D(D_21), .E(n6268), .C(wclk), .QN(n3579) );
  DFE1 \mem_reg_106][20  ( .D(D_20), .E(n6268), .C(wclk), .QN(n3580) );
  DFE1 \mem_reg_106][19  ( .D(D_19), .E(n6268), .C(wclk), .QN(n3581) );
  DFE1 \mem_reg_106][18  ( .D(D_18), .E(n6268), .C(wclk), .QN(n3582) );
  DFE1 \mem_reg_106][17  ( .D(D_17), .E(n6268), .C(wclk), .QN(n3583) );
  DFE1 \mem_reg_106][16  ( .D(D_16), .E(n6268), .C(wclk), .QN(n3584) );
  DFE1 \mem_reg_106][15  ( .D(D_15), .E(n6268), .C(wclk), .QN(n3585) );
  DFE1 \mem_reg_106][14  ( .D(D_14), .E(n6268), .C(wclk), .QN(n3586) );
  DFE1 \mem_reg_106][13  ( .D(D_13), .E(n6268), .C(wclk), .QN(n3587) );
  DFE1 \mem_reg_106][12  ( .D(D_12), .E(n6268), .C(wclk), .QN(n3588) );
  DFE1 \mem_reg_106][11  ( .D(D_11), .E(n6268), .C(wclk), .QN(n3589) );
  DFE1 \mem_reg_106][10  ( .D(D_10), .E(n6268), .C(wclk), .QN(n3590) );
  DFE1 \mem_reg_106][9  ( .D(D_9), .E(n6268), .C(wclk), .QN(n3591) );
  DFE1 \mem_reg_106][8  ( .D(D_8), .E(n6268), .C(wclk), .QN(n3592) );
  DFE1 \mem_reg_106][7  ( .D(D_7), .E(n6268), .C(wclk), .QN(n3593) );
  DFE1 \mem_reg_106][6  ( .D(D_6), .E(n6268), .C(wclk), .QN(n3594) );
  DFE1 \mem_reg_106][5  ( .D(D_5), .E(n6268), .C(wclk), .QN(n3595) );
  DFE1 \mem_reg_106][4  ( .D(D_4), .E(n6268), .C(wclk), .QN(n3596) );
  DFE1 \mem_reg_106][3  ( .D(D_3), .E(n6268), .C(wclk), .QN(n3597) );
  DFE1 \mem_reg_106][2  ( .D(D_2), .E(n6268), .C(wclk), .QN(n3598) );
  DFE1 \mem_reg_106][1  ( .D(D_1), .E(n6268), .C(wclk), .QN(n3599) );
  DFE1 \mem_reg_106][0  ( .D(D_0), .E(n6268), .C(wclk), .QN(n3600) );
  DFE1 \mem_reg_105][23  ( .D(D_23), .E(n6267), .C(wclk), .QN(n3601) );
  DFE1 \mem_reg_105][22  ( .D(D_22), .E(n6267), .C(wclk), .QN(n3602) );
  DFE1 \mem_reg_105][21  ( .D(D_21), .E(n6267), .C(wclk), .QN(n3603) );
  DFE1 \mem_reg_105][20  ( .D(D_20), .E(n6267), .C(wclk), .QN(n3604) );
  DFE1 \mem_reg_105][19  ( .D(D_19), .E(n6267), .C(wclk), .QN(n3605) );
  DFE1 \mem_reg_105][18  ( .D(D_18), .E(n6267), .C(wclk), .QN(n3606) );
  DFE1 \mem_reg_105][17  ( .D(D_17), .E(n6267), .C(wclk), .QN(n3607) );
  DFE1 \mem_reg_105][16  ( .D(D_16), .E(n6267), .C(wclk), .QN(n3608) );
  DFE1 \mem_reg_105][15  ( .D(D_15), .E(n6267), .C(wclk), .QN(n3609) );
  DFE1 \mem_reg_105][14  ( .D(D_14), .E(n6267), .C(wclk), .QN(n3610) );
  DFE1 \mem_reg_105][13  ( .D(D_13), .E(n6267), .C(wclk), .QN(n3611) );
  DFE1 \mem_reg_105][12  ( .D(D_12), .E(n6267), .C(wclk), .QN(n3612) );
  DFE1 \mem_reg_105][11  ( .D(D_11), .E(n6267), .C(wclk), .QN(n3613) );
  DFE1 \mem_reg_105][10  ( .D(D_10), .E(n6267), .C(wclk), .QN(n3614) );
  DFE1 \mem_reg_105][9  ( .D(D_9), .E(n6267), .C(wclk), .QN(n3615) );
  DFE1 \mem_reg_105][8  ( .D(D_8), .E(n6267), .C(wclk), .QN(n3616) );
  DFE1 \mem_reg_105][7  ( .D(D_7), .E(n6267), .C(wclk), .QN(n3617) );
  DFE1 \mem_reg_105][6  ( .D(D_6), .E(n6267), .C(wclk), .QN(n3618) );
  DFE1 \mem_reg_105][5  ( .D(D_5), .E(n6267), .C(wclk), .QN(n3619) );
  DFE1 \mem_reg_105][4  ( .D(D_4), .E(n6267), .C(wclk), .QN(n3620) );
  DFE1 \mem_reg_105][3  ( .D(D_3), .E(n6267), .C(wclk), .QN(n3621) );
  DFE1 \mem_reg_105][2  ( .D(D_2), .E(n6267), .C(wclk), .QN(n3622) );
  DFE1 \mem_reg_105][1  ( .D(D_1), .E(n6267), .C(wclk), .QN(n3623) );
  DFE1 \mem_reg_105][0  ( .D(D_0), .E(n6267), .C(wclk), .QN(n3624) );
  DFE1 \mem_reg_104][23  ( .D(D_23), .E(n6266), .C(wclk), .QN(n3625) );
  DFE1 \mem_reg_104][22  ( .D(D_22), .E(n6266), .C(wclk), .QN(n3626) );
  DFE1 \mem_reg_104][21  ( .D(D_21), .E(n6266), .C(wclk), .QN(n3627) );
  DFE1 \mem_reg_104][20  ( .D(D_20), .E(n6266), .C(wclk), .QN(n3628) );
  DFE1 \mem_reg_104][19  ( .D(D_19), .E(n6266), .C(wclk), .QN(n3629) );
  DFE1 \mem_reg_104][18  ( .D(D_18), .E(n6266), .C(wclk), .QN(n3630) );
  DFE1 \mem_reg_104][17  ( .D(D_17), .E(n6266), .C(wclk), .QN(n3631) );
  DFE1 \mem_reg_104][16  ( .D(D_16), .E(n6266), .C(wclk), .QN(n3632) );
  DFE1 \mem_reg_104][15  ( .D(D_15), .E(n6266), .C(wclk), .QN(n3633) );
  DFE1 \mem_reg_104][14  ( .D(D_14), .E(n6266), .C(wclk), .QN(n3634) );
  DFE1 \mem_reg_104][13  ( .D(D_13), .E(n6266), .C(wclk), .QN(n3635) );
  DFE1 \mem_reg_104][12  ( .D(D_12), .E(n6266), .C(wclk), .QN(n3636) );
  DFE1 \mem_reg_104][11  ( .D(D_11), .E(n6266), .C(wclk), .QN(n3637) );
  DFE1 \mem_reg_104][10  ( .D(D_10), .E(n6266), .C(wclk), .QN(n3638) );
  DFE1 \mem_reg_104][9  ( .D(D_9), .E(n6266), .C(wclk), .QN(n3639) );
  DFE1 \mem_reg_104][8  ( .D(D_8), .E(n6266), .C(wclk), .QN(n3640) );
  DFE1 \mem_reg_104][7  ( .D(D_7), .E(n6266), .C(wclk), .QN(n3641) );
  DFE1 \mem_reg_104][6  ( .D(D_6), .E(n6266), .C(wclk), .QN(n3642) );
  DFE1 \mem_reg_104][5  ( .D(D_5), .E(n6266), .C(wclk), .QN(n3643) );
  DFE1 \mem_reg_104][4  ( .D(D_4), .E(n6266), .C(wclk), .QN(n3644) );
  DFE1 \mem_reg_104][3  ( .D(D_3), .E(n6266), .C(wclk), .QN(n3645) );
  DFE1 \mem_reg_104][2  ( .D(D_2), .E(n6266), .C(wclk), .QN(n3646) );
  DFE1 \mem_reg_104][1  ( .D(D_1), .E(n6266), .C(wclk), .QN(n3647) );
  DFE1 \mem_reg_104][0  ( .D(D_0), .E(n6266), .C(wclk), .QN(n3648) );
  DFE1 \mem_reg_103][23  ( .D(D_23), .E(n6264), .C(wclk), .QN(n3649) );
  DFE1 \mem_reg_103][22  ( .D(D_22), .E(n6264), .C(wclk), .QN(n3650) );
  DFE1 \mem_reg_103][21  ( .D(D_21), .E(n6264), .C(wclk), .QN(n3651) );
  DFE1 \mem_reg_103][20  ( .D(D_20), .E(n6264), .C(wclk), .QN(n3652) );
  DFE1 \mem_reg_103][19  ( .D(D_19), .E(n6264), .C(wclk), .QN(n3653) );
  DFE1 \mem_reg_103][18  ( .D(D_18), .E(n6264), .C(wclk), .QN(n3654) );
  DFE1 \mem_reg_103][17  ( .D(D_17), .E(n6264), .C(wclk), .QN(n3655) );
  DFE1 \mem_reg_103][16  ( .D(D_16), .E(n6264), .C(wclk), .QN(n3656) );
  DFE1 \mem_reg_103][15  ( .D(D_15), .E(n6264), .C(wclk), .QN(n3657) );
  DFE1 \mem_reg_103][14  ( .D(D_14), .E(n6264), .C(wclk), .QN(n3658) );
  DFE1 \mem_reg_103][13  ( .D(D_13), .E(n6264), .C(wclk), .QN(n3659) );
  DFE1 \mem_reg_103][12  ( .D(D_12), .E(n6264), .C(wclk), .QN(n3660) );
  DFE1 \mem_reg_103][11  ( .D(D_11), .E(n6264), .C(wclk), .QN(n3661) );
  DFE1 \mem_reg_103][10  ( .D(D_10), .E(n6264), .C(wclk), .QN(n3662) );
  DFE1 \mem_reg_103][9  ( .D(D_9), .E(n6264), .C(wclk), .QN(n3663) );
  DFE1 \mem_reg_103][8  ( .D(D_8), .E(n6264), .C(wclk), .QN(n3664) );
  DFE1 \mem_reg_103][7  ( .D(D_7), .E(n6264), .C(wclk), .QN(n3665) );
  DFE1 \mem_reg_103][6  ( .D(D_6), .E(n6264), .C(wclk), .QN(n3666) );
  DFE1 \mem_reg_103][5  ( .D(D_5), .E(n6264), .C(wclk), .QN(n3667) );
  DFE1 \mem_reg_103][4  ( .D(D_4), .E(n6264), .C(wclk), .QN(n3668) );
  DFE1 \mem_reg_103][3  ( .D(D_3), .E(n6264), .C(wclk), .QN(n3669) );
  DFE1 \mem_reg_103][2  ( .D(D_2), .E(n6264), .C(wclk), .QN(n3670) );
  DFE1 \mem_reg_103][1  ( .D(D_1), .E(n6264), .C(wclk), .QN(n3671) );
  DFE1 \mem_reg_103][0  ( .D(D_0), .E(n6264), .C(wclk), .QN(n3672) );
  DFE1 \mem_reg_102][23  ( .D(D_23), .E(n6263), .C(wclk), .QN(n3673) );
  DFE1 \mem_reg_102][22  ( .D(D_22), .E(n6263), .C(wclk), .QN(n3674) );
  DFE1 \mem_reg_102][21  ( .D(D_21), .E(n6263), .C(wclk), .QN(n3675) );
  DFE1 \mem_reg_102][20  ( .D(D_20), .E(n6263), .C(wclk), .QN(n3676) );
  DFE1 \mem_reg_102][19  ( .D(D_19), .E(n6263), .C(wclk), .QN(n3677) );
  DFE1 \mem_reg_102][18  ( .D(D_18), .E(n6263), .C(wclk), .QN(n3678) );
  DFE1 \mem_reg_102][17  ( .D(D_17), .E(n6263), .C(wclk), .QN(n3679) );
  DFE1 \mem_reg_102][16  ( .D(D_16), .E(n6263), .C(wclk), .QN(n3680) );
  DFE1 \mem_reg_102][15  ( .D(D_15), .E(n6263), .C(wclk), .QN(n3681) );
  DFE1 \mem_reg_102][14  ( .D(D_14), .E(n6263), .C(wclk), .QN(n3682) );
  DFE1 \mem_reg_102][13  ( .D(D_13), .E(n6263), .C(wclk), .QN(n3683) );
  DFE1 \mem_reg_102][12  ( .D(D_12), .E(n6263), .C(wclk), .QN(n3684) );
  DFE1 \mem_reg_102][11  ( .D(D_11), .E(n6263), .C(wclk), .QN(n3685) );
  DFE1 \mem_reg_102][10  ( .D(D_10), .E(n6263), .C(wclk), .QN(n3686) );
  DFE1 \mem_reg_102][9  ( .D(D_9), .E(n6263), .C(wclk), .QN(n3687) );
  DFE1 \mem_reg_102][8  ( .D(D_8), .E(n6263), .C(wclk), .QN(n3688) );
  DFE1 \mem_reg_102][7  ( .D(D_7), .E(n6263), .C(wclk), .QN(n3689) );
  DFE1 \mem_reg_102][6  ( .D(D_6), .E(n6263), .C(wclk), .QN(n3690) );
  DFE1 \mem_reg_102][5  ( .D(D_5), .E(n6263), .C(wclk), .QN(n3691) );
  DFE1 \mem_reg_102][4  ( .D(D_4), .E(n6263), .C(wclk), .QN(n3692) );
  DFE1 \mem_reg_102][3  ( .D(D_3), .E(n6263), .C(wclk), .QN(n3693) );
  DFE1 \mem_reg_102][2  ( .D(D_2), .E(n6263), .C(wclk), .QN(n3694) );
  DFE1 \mem_reg_102][1  ( .D(D_1), .E(n6263), .C(wclk), .QN(n3695) );
  DFE1 \mem_reg_102][0  ( .D(D_0), .E(n6263), .C(wclk), .QN(n3696) );
  DFE1 \mem_reg_101][23  ( .D(D_23), .E(n6262), .C(wclk), .QN(n3697) );
  DFE1 \mem_reg_101][22  ( .D(D_22), .E(n6262), .C(wclk), .QN(n3698) );
  DFE1 \mem_reg_101][21  ( .D(D_21), .E(n6262), .C(wclk), .QN(n3699) );
  DFE1 \mem_reg_101][20  ( .D(D_20), .E(n6262), .C(wclk), .QN(n3700) );
  DFE1 \mem_reg_101][19  ( .D(D_19), .E(n6262), .C(wclk), .QN(n3701) );
  DFE1 \mem_reg_101][18  ( .D(D_18), .E(n6262), .C(wclk), .QN(n3702) );
  DFE1 \mem_reg_101][17  ( .D(D_17), .E(n6262), .C(wclk), .QN(n3703) );
  DFE1 \mem_reg_101][16  ( .D(D_16), .E(n6262), .C(wclk), .QN(n3704) );
  DFE1 \mem_reg_101][15  ( .D(D_15), .E(n6262), .C(wclk), .QN(n3705) );
  DFE1 \mem_reg_101][14  ( .D(D_14), .E(n6262), .C(wclk), .QN(n3706) );
  DFE1 \mem_reg_101][13  ( .D(D_13), .E(n6262), .C(wclk), .QN(n3707) );
  DFE1 \mem_reg_101][12  ( .D(D_12), .E(n6262), .C(wclk), .QN(n3708) );
  DFE1 \mem_reg_101][11  ( .D(D_11), .E(n6262), .C(wclk), .QN(n3709) );
  DFE1 \mem_reg_101][10  ( .D(D_10), .E(n6262), .C(wclk), .QN(n3710) );
  DFE1 \mem_reg_101][9  ( .D(D_9), .E(n6262), .C(wclk), .QN(n3711) );
  DFE1 \mem_reg_101][8  ( .D(D_8), .E(n6262), .C(wclk), .QN(n3712) );
  DFE1 \mem_reg_101][7  ( .D(D_7), .E(n6262), .C(wclk), .QN(n3713) );
  DFE1 \mem_reg_101][6  ( .D(D_6), .E(n6262), .C(wclk), .QN(n3714) );
  DFE1 \mem_reg_101][5  ( .D(D_5), .E(n6262), .C(wclk), .QN(n3715) );
  DFE1 \mem_reg_101][4  ( .D(D_4), .E(n6262), .C(wclk), .QN(n3716) );
  DFE1 \mem_reg_101][3  ( .D(D_3), .E(n6262), .C(wclk), .QN(n3717) );
  DFE1 \mem_reg_101][2  ( .D(D_2), .E(n6262), .C(wclk), .QN(n3718) );
  DFE1 \mem_reg_101][1  ( .D(D_1), .E(n6262), .C(wclk), .QN(n3719) );
  DFE1 \mem_reg_101][0  ( .D(D_0), .E(n6262), .C(wclk), .QN(n3720) );
  DFE1 \mem_reg_100][23  ( .D(D_23), .E(n6261), .C(wclk), .QN(n3721) );
  DFE1 \mem_reg_100][22  ( .D(D_22), .E(n6261), .C(wclk), .QN(n3722) );
  DFE1 \mem_reg_100][21  ( .D(D_21), .E(n6261), .C(wclk), .QN(n3723) );
  DFE1 \mem_reg_100][20  ( .D(D_20), .E(n6261), .C(wclk), .QN(n3724) );
  DFE1 \mem_reg_100][19  ( .D(D_19), .E(n6261), .C(wclk), .QN(n3725) );
  DFE1 \mem_reg_100][18  ( .D(D_18), .E(n6261), .C(wclk), .QN(n3726) );
  DFE1 \mem_reg_100][17  ( .D(D_17), .E(n6261), .C(wclk), .QN(n3727) );
  DFE1 \mem_reg_100][16  ( .D(D_16), .E(n6261), .C(wclk), .QN(n3728) );
  DFE1 \mem_reg_100][15  ( .D(D_15), .E(n6261), .C(wclk), .QN(n3729) );
  DFE1 \mem_reg_100][14  ( .D(D_14), .E(n6261), .C(wclk), .QN(n3730) );
  DFE1 \mem_reg_100][13  ( .D(D_13), .E(n6261), .C(wclk), .QN(n3731) );
  DFE1 \mem_reg_100][12  ( .D(D_12), .E(n6261), .C(wclk), .QN(n3732) );
  DFE1 \mem_reg_100][11  ( .D(D_11), .E(n6261), .C(wclk), .QN(n3733) );
  DFE1 \mem_reg_100][10  ( .D(D_10), .E(n6261), .C(wclk), .QN(n3734) );
  DFE1 \mem_reg_100][9  ( .D(D_9), .E(n6261), .C(wclk), .QN(n3735) );
  DFE1 \mem_reg_100][8  ( .D(D_8), .E(n6261), .C(wclk), .QN(n3736) );
  DFE1 \mem_reg_100][7  ( .D(D_7), .E(n6261), .C(wclk), .QN(n3737) );
  DFE1 \mem_reg_100][6  ( .D(D_6), .E(n6261), .C(wclk), .QN(n3738) );
  DFE1 \mem_reg_100][5  ( .D(D_5), .E(n6261), .C(wclk), .QN(n3739) );
  DFE1 \mem_reg_100][4  ( .D(D_4), .E(n6261), .C(wclk), .QN(n3740) );
  DFE1 \mem_reg_100][3  ( .D(D_3), .E(n6261), .C(wclk), .QN(n3741) );
  DFE1 \mem_reg_100][2  ( .D(D_2), .E(n6261), .C(wclk), .QN(n3742) );
  DFE1 \mem_reg_100][1  ( .D(D_1), .E(n6261), .C(wclk), .QN(n3743) );
  DFE1 \mem_reg_100][0  ( .D(D_0), .E(n6261), .C(wclk), .QN(n3744) );
  DFE1 \mem_reg_99][23  ( .D(D_23), .E(n6260), .C(wclk), .QN(n3745) );
  DFE1 \mem_reg_99][22  ( .D(D_22), .E(n6260), .C(wclk), .QN(n3746) );
  DFE1 \mem_reg_99][21  ( .D(D_21), .E(n6260), .C(wclk), .QN(n3747) );
  DFE1 \mem_reg_99][20  ( .D(D_20), .E(n6260), .C(wclk), .QN(n3748) );
  DFE1 \mem_reg_99][19  ( .D(D_19), .E(n6260), .C(wclk), .QN(n3749) );
  DFE1 \mem_reg_99][18  ( .D(D_18), .E(n6260), .C(wclk), .QN(n3750) );
  DFE1 \mem_reg_99][17  ( .D(D_17), .E(n6260), .C(wclk), .QN(n3751) );
  DFE1 \mem_reg_99][16  ( .D(D_16), .E(n6260), .C(wclk), .QN(n3752) );
  DFE1 \mem_reg_99][15  ( .D(D_15), .E(n6260), .C(wclk), .QN(n3753) );
  DFE1 \mem_reg_99][14  ( .D(D_14), .E(n6260), .C(wclk), .QN(n3754) );
  DFE1 \mem_reg_99][13  ( .D(D_13), .E(n6260), .C(wclk), .QN(n3755) );
  DFE1 \mem_reg_99][12  ( .D(D_12), .E(n6260), .C(wclk), .QN(n3756) );
  DFE1 \mem_reg_99][11  ( .D(D_11), .E(n6260), .C(wclk), .QN(n3757) );
  DFE1 \mem_reg_99][10  ( .D(D_10), .E(n6260), .C(wclk), .QN(n3758) );
  DFE1 \mem_reg_99][9  ( .D(D_9), .E(n6260), .C(wclk), .QN(n3759) );
  DFE1 \mem_reg_99][8  ( .D(D_8), .E(n6260), .C(wclk), .QN(n3760) );
  DFE1 \mem_reg_99][7  ( .D(D_7), .E(n6260), .C(wclk), .QN(n3761) );
  DFE1 \mem_reg_99][6  ( .D(D_6), .E(n6260), .C(wclk), .QN(n3762) );
  DFE1 \mem_reg_99][5  ( .D(D_5), .E(n6260), .C(wclk), .QN(n3763) );
  DFE1 \mem_reg_99][4  ( .D(D_4), .E(n6260), .C(wclk), .QN(n3764) );
  DFE1 \mem_reg_99][3  ( .D(D_3), .E(n6260), .C(wclk), .QN(n3765) );
  DFE1 \mem_reg_99][2  ( .D(D_2), .E(n6260), .C(wclk), .QN(n3766) );
  DFE1 \mem_reg_99][1  ( .D(D_1), .E(n6260), .C(wclk), .QN(n3767) );
  DFE1 \mem_reg_99][0  ( .D(D_0), .E(n6260), .C(wclk), .QN(n3768) );
  DFE1 \mem_reg_98][23  ( .D(D_23), .E(n6259), .C(wclk), .QN(n3769) );
  DFE1 \mem_reg_98][22  ( .D(D_22), .E(n6259), .C(wclk), .QN(n3770) );
  DFE1 \mem_reg_98][21  ( .D(D_21), .E(n6259), .C(wclk), .QN(n3771) );
  DFE1 \mem_reg_98][20  ( .D(D_20), .E(n6259), .C(wclk), .QN(n3772) );
  DFE1 \mem_reg_98][19  ( .D(D_19), .E(n6259), .C(wclk), .QN(n3773) );
  DFE1 \mem_reg_98][18  ( .D(D_18), .E(n6259), .C(wclk), .QN(n3774) );
  DFE1 \mem_reg_98][17  ( .D(D_17), .E(n6259), .C(wclk), .QN(n3775) );
  DFE1 \mem_reg_98][16  ( .D(D_16), .E(n6259), .C(wclk), .QN(n3776) );
  DFE1 \mem_reg_98][15  ( .D(D_15), .E(n6259), .C(wclk), .QN(n3777) );
  DFE1 \mem_reg_98][14  ( .D(D_14), .E(n6259), .C(wclk), .QN(n3778) );
  DFE1 \mem_reg_98][13  ( .D(D_13), .E(n6259), .C(wclk), .QN(n3779) );
  DFE1 \mem_reg_98][12  ( .D(D_12), .E(n6259), .C(wclk), .QN(n3780) );
  DFE1 \mem_reg_98][11  ( .D(D_11), .E(n6259), .C(wclk), .QN(n3781) );
  DFE1 \mem_reg_98][10  ( .D(D_10), .E(n6259), .C(wclk), .QN(n3782) );
  DFE1 \mem_reg_98][9  ( .D(D_9), .E(n6259), .C(wclk), .QN(n3783) );
  DFE1 \mem_reg_98][8  ( .D(D_8), .E(n6259), .C(wclk), .QN(n3784) );
  DFE1 \mem_reg_98][7  ( .D(D_7), .E(n6259), .C(wclk), .QN(n3785) );
  DFE1 \mem_reg_98][6  ( .D(D_6), .E(n6259), .C(wclk), .QN(n3786) );
  DFE1 \mem_reg_98][5  ( .D(D_5), .E(n6259), .C(wclk), .QN(n3787) );
  DFE1 \mem_reg_98][4  ( .D(D_4), .E(n6259), .C(wclk), .QN(n3788) );
  DFE1 \mem_reg_98][3  ( .D(D_3), .E(n6259), .C(wclk), .QN(n3789) );
  DFE1 \mem_reg_98][2  ( .D(D_2), .E(n6259), .C(wclk), .QN(n3790) );
  DFE1 \mem_reg_98][1  ( .D(D_1), .E(n6259), .C(wclk), .QN(n3791) );
  DFE1 \mem_reg_98][0  ( .D(D_0), .E(n6259), .C(wclk), .QN(n3792) );
  DFE1 \mem_reg_97][23  ( .D(D_23), .E(n6258), .C(wclk), .QN(n3793) );
  DFE1 \mem_reg_97][22  ( .D(D_22), .E(n6258), .C(wclk), .QN(n3794) );
  DFE1 \mem_reg_97][21  ( .D(D_21), .E(n6258), .C(wclk), .QN(n3795) );
  DFE1 \mem_reg_97][20  ( .D(D_20), .E(n6258), .C(wclk), .QN(n3796) );
  DFE1 \mem_reg_97][19  ( .D(D_19), .E(n6258), .C(wclk), .QN(n3797) );
  DFE1 \mem_reg_97][18  ( .D(D_18), .E(n6258), .C(wclk), .QN(n3798) );
  DFE1 \mem_reg_97][17  ( .D(D_17), .E(n6258), .C(wclk), .QN(n3799) );
  DFE1 \mem_reg_97][16  ( .D(D_16), .E(n6258), .C(wclk), .QN(n3800) );
  DFE1 \mem_reg_97][15  ( .D(D_15), .E(n6258), .C(wclk), .QN(n3801) );
  DFE1 \mem_reg_97][14  ( .D(D_14), .E(n6258), .C(wclk), .QN(n3802) );
  DFE1 \mem_reg_97][13  ( .D(D_13), .E(n6258), .C(wclk), .QN(n3803) );
  DFE1 \mem_reg_97][12  ( .D(D_12), .E(n6258), .C(wclk), .QN(n3804) );
  DFE1 \mem_reg_97][11  ( .D(D_11), .E(n6258), .C(wclk), .QN(n3805) );
  DFE1 \mem_reg_97][10  ( .D(D_10), .E(n6258), .C(wclk), .QN(n3806) );
  DFE1 \mem_reg_97][9  ( .D(D_9), .E(n6258), .C(wclk), .QN(n3807) );
  DFE1 \mem_reg_97][8  ( .D(D_8), .E(n6258), .C(wclk), .QN(n3808) );
  DFE1 \mem_reg_97][7  ( .D(D_7), .E(n6258), .C(wclk), .QN(n3809) );
  DFE1 \mem_reg_97][6  ( .D(D_6), .E(n6258), .C(wclk), .QN(n3810) );
  DFE1 \mem_reg_97][5  ( .D(D_5), .E(n6258), .C(wclk), .QN(n3811) );
  DFE1 \mem_reg_97][4  ( .D(D_4), .E(n6258), .C(wclk), .QN(n3812) );
  DFE1 \mem_reg_97][3  ( .D(D_3), .E(n6258), .C(wclk), .QN(n3813) );
  DFE1 \mem_reg_97][2  ( .D(D_2), .E(n6258), .C(wclk), .QN(n3814) );
  DFE1 \mem_reg_97][1  ( .D(D_1), .E(n6258), .C(wclk), .QN(n3815) );
  DFE1 \mem_reg_97][0  ( .D(D_0), .E(n6258), .C(wclk), .QN(n3816) );
  DFE1 \mem_reg_96][23  ( .D(D_23), .E(n6256), .C(wclk), .QN(n3817) );
  DFE1 \mem_reg_96][22  ( .D(D_22), .E(n6256), .C(wclk), .QN(n3818) );
  DFE1 \mem_reg_96][21  ( .D(D_21), .E(n6256), .C(wclk), .QN(n3819) );
  DFE1 \mem_reg_96][20  ( .D(D_20), .E(n6256), .C(wclk), .QN(n3820) );
  DFE1 \mem_reg_96][19  ( .D(D_19), .E(n6256), .C(wclk), .QN(n3821) );
  DFE1 \mem_reg_96][18  ( .D(D_18), .E(n6256), .C(wclk), .QN(n3822) );
  DFE1 \mem_reg_96][17  ( .D(D_17), .E(n6256), .C(wclk), .QN(n3823) );
  DFE1 \mem_reg_96][16  ( .D(D_16), .E(n6256), .C(wclk), .QN(n3824) );
  DFE1 \mem_reg_96][15  ( .D(D_15), .E(n6256), .C(wclk), .QN(n3825) );
  DFE1 \mem_reg_96][14  ( .D(D_14), .E(n6256), .C(wclk), .QN(n3826) );
  DFE1 \mem_reg_96][13  ( .D(D_13), .E(n6256), .C(wclk), .QN(n3827) );
  DFE1 \mem_reg_96][12  ( .D(D_12), .E(n6256), .C(wclk), .QN(n3828) );
  DFE1 \mem_reg_96][11  ( .D(D_11), .E(n6256), .C(wclk), .QN(n3829) );
  DFE1 \mem_reg_96][10  ( .D(D_10), .E(n6256), .C(wclk), .QN(n3830) );
  DFE1 \mem_reg_96][9  ( .D(D_9), .E(n6256), .C(wclk), .QN(n3831) );
  DFE1 \mem_reg_96][8  ( .D(D_8), .E(n6256), .C(wclk), .QN(n3832) );
  DFE1 \mem_reg_96][7  ( .D(D_7), .E(n6256), .C(wclk), .QN(n3833) );
  DFE1 \mem_reg_96][6  ( .D(D_6), .E(n6256), .C(wclk), .QN(n3834) );
  DFE1 \mem_reg_96][5  ( .D(D_5), .E(n6256), .C(wclk), .QN(n3835) );
  DFE1 \mem_reg_96][4  ( .D(D_4), .E(n6256), .C(wclk), .QN(n3836) );
  DFE1 \mem_reg_96][3  ( .D(D_3), .E(n6256), .C(wclk), .QN(n3837) );
  DFE1 \mem_reg_96][2  ( .D(D_2), .E(n6256), .C(wclk), .QN(n3838) );
  DFE1 \mem_reg_96][1  ( .D(D_1), .E(n6256), .C(wclk), .QN(n3839) );
  DFE1 \mem_reg_96][0  ( .D(D_0), .E(n6256), .C(wclk), .QN(n3840) );
  DFE1 \mem_reg_95][23  ( .D(D_23), .E(n6254), .C(wclk), .QN(n3841) );
  DFE1 \mem_reg_95][22  ( .D(D_22), .E(n6254), .C(wclk), .QN(n3842) );
  DFE1 \mem_reg_95][21  ( .D(D_21), .E(n6254), .C(wclk), .QN(n3843) );
  DFE1 \mem_reg_95][20  ( .D(D_20), .E(n6254), .C(wclk), .QN(n3844) );
  DFE1 \mem_reg_95][19  ( .D(D_19), .E(n6254), .C(wclk), .QN(n3845) );
  DFE1 \mem_reg_95][18  ( .D(D_18), .E(n6254), .C(wclk), .QN(n3846) );
  DFE1 \mem_reg_95][17  ( .D(D_17), .E(n6254), .C(wclk), .QN(n3847) );
  DFE1 \mem_reg_95][16  ( .D(D_16), .E(n6254), .C(wclk), .QN(n3848) );
  DFE1 \mem_reg_95][15  ( .D(D_15), .E(n6254), .C(wclk), .QN(n3849) );
  DFE1 \mem_reg_95][14  ( .D(D_14), .E(n6254), .C(wclk), .QN(n3850) );
  DFE1 \mem_reg_95][13  ( .D(D_13), .E(n6254), .C(wclk), .QN(n3851) );
  DFE1 \mem_reg_95][12  ( .D(D_12), .E(n6254), .C(wclk), .QN(n3852) );
  DFE1 \mem_reg_95][11  ( .D(D_11), .E(n6254), .C(wclk), .QN(n3853) );
  DFE1 \mem_reg_95][10  ( .D(D_10), .E(n6254), .C(wclk), .QN(n3854) );
  DFE1 \mem_reg_95][9  ( .D(D_9), .E(n6254), .C(wclk), .QN(n3855) );
  DFE1 \mem_reg_95][8  ( .D(D_8), .E(n6254), .C(wclk), .QN(n3856) );
  DFE1 \mem_reg_95][7  ( .D(D_7), .E(n6254), .C(wclk), .QN(n3857) );
  DFE1 \mem_reg_95][6  ( .D(D_6), .E(n6254), .C(wclk), .QN(n3858) );
  DFE1 \mem_reg_95][5  ( .D(D_5), .E(n6254), .C(wclk), .QN(n3859) );
  DFE1 \mem_reg_95][4  ( .D(D_4), .E(n6254), .C(wclk), .QN(n3860) );
  DFE1 \mem_reg_95][3  ( .D(D_3), .E(n6254), .C(wclk), .QN(n3861) );
  DFE1 \mem_reg_95][2  ( .D(D_2), .E(n6254), .C(wclk), .QN(n3862) );
  DFE1 \mem_reg_95][1  ( .D(D_1), .E(n6254), .C(wclk), .QN(n3863) );
  DFE1 \mem_reg_95][0  ( .D(D_0), .E(n6254), .C(wclk), .QN(n3864) );
  DFE1 \mem_reg_94][23  ( .D(D_23), .E(n6253), .C(wclk), .QN(n3865) );
  DFE1 \mem_reg_94][22  ( .D(D_22), .E(n6253), .C(wclk), .QN(n3866) );
  DFE1 \mem_reg_94][21  ( .D(D_21), .E(n6253), .C(wclk), .QN(n3867) );
  DFE1 \mem_reg_94][20  ( .D(D_20), .E(n6253), .C(wclk), .QN(n3868) );
  DFE1 \mem_reg_94][19  ( .D(D_19), .E(n6253), .C(wclk), .QN(n3869) );
  DFE1 \mem_reg_94][18  ( .D(D_18), .E(n6253), .C(wclk), .QN(n3870) );
  DFE1 \mem_reg_94][17  ( .D(D_17), .E(n6253), .C(wclk), .QN(n3871) );
  DFE1 \mem_reg_94][16  ( .D(D_16), .E(n6253), .C(wclk), .QN(n3872) );
  DFE1 \mem_reg_94][15  ( .D(D_15), .E(n6253), .C(wclk), .QN(n3873) );
  DFE1 \mem_reg_94][14  ( .D(D_14), .E(n6253), .C(wclk), .QN(n3874) );
  DFE1 \mem_reg_94][13  ( .D(D_13), .E(n6253), .C(wclk), .QN(n3875) );
  DFE1 \mem_reg_94][12  ( .D(D_12), .E(n6253), .C(wclk), .QN(n3876) );
  DFE1 \mem_reg_94][11  ( .D(D_11), .E(n6253), .C(wclk), .QN(n3877) );
  DFE1 \mem_reg_94][10  ( .D(D_10), .E(n6253), .C(wclk), .QN(n3878) );
  DFE1 \mem_reg_94][9  ( .D(D_9), .E(n6253), .C(wclk), .QN(n3879) );
  DFE1 \mem_reg_94][8  ( .D(D_8), .E(n6253), .C(wclk), .QN(n3880) );
  DFE1 \mem_reg_94][7  ( .D(D_7), .E(n6253), .C(wclk), .QN(n3881) );
  DFE1 \mem_reg_94][6  ( .D(D_6), .E(n6253), .C(wclk), .QN(n3882) );
  DFE1 \mem_reg_94][5  ( .D(D_5), .E(n6253), .C(wclk), .QN(n3883) );
  DFE1 \mem_reg_94][4  ( .D(D_4), .E(n6253), .C(wclk), .QN(n3884) );
  DFE1 \mem_reg_94][3  ( .D(D_3), .E(n6253), .C(wclk), .QN(n3885) );
  DFE1 \mem_reg_94][2  ( .D(D_2), .E(n6253), .C(wclk), .QN(n3886) );
  DFE1 \mem_reg_94][1  ( .D(D_1), .E(n6253), .C(wclk), .QN(n3887) );
  DFE1 \mem_reg_94][0  ( .D(D_0), .E(n6253), .C(wclk), .QN(n3888) );
  DFE1 \mem_reg_93][23  ( .D(D_23), .E(n6251), .C(wclk), .QN(n3889) );
  DFE1 \mem_reg_93][22  ( .D(D_22), .E(n6251), .C(wclk), .QN(n3890) );
  DFE1 \mem_reg_93][21  ( .D(D_21), .E(n6251), .C(wclk), .QN(n3891) );
  DFE1 \mem_reg_93][20  ( .D(D_20), .E(n6251), .C(wclk), .QN(n3892) );
  DFE1 \mem_reg_93][19  ( .D(D_19), .E(n6251), .C(wclk), .QN(n3893) );
  DFE1 \mem_reg_93][18  ( .D(D_18), .E(n6251), .C(wclk), .QN(n3894) );
  DFE1 \mem_reg_93][17  ( .D(D_17), .E(n6251), .C(wclk), .QN(n3895) );
  DFE1 \mem_reg_93][16  ( .D(D_16), .E(n6251), .C(wclk), .QN(n3896) );
  DFE1 \mem_reg_93][15  ( .D(D_15), .E(n6251), .C(wclk), .QN(n3897) );
  DFE1 \mem_reg_93][14  ( .D(D_14), .E(n6251), .C(wclk), .QN(n3898) );
  DFE1 \mem_reg_93][13  ( .D(D_13), .E(n6251), .C(wclk), .QN(n3899) );
  DFE1 \mem_reg_93][12  ( .D(D_12), .E(n6251), .C(wclk), .QN(n3900) );
  DFE1 \mem_reg_93][11  ( .D(D_11), .E(n6251), .C(wclk), .QN(n3901) );
  DFE1 \mem_reg_93][10  ( .D(D_10), .E(n6251), .C(wclk), .QN(n3902) );
  DFE1 \mem_reg_93][9  ( .D(D_9), .E(n6251), .C(wclk), .QN(n3903) );
  DFE1 \mem_reg_93][8  ( .D(D_8), .E(n6251), .C(wclk), .QN(n3904) );
  DFE1 \mem_reg_93][7  ( .D(D_7), .E(n6251), .C(wclk), .QN(n3905) );
  DFE1 \mem_reg_93][6  ( .D(D_6), .E(n6251), .C(wclk), .QN(n3906) );
  DFE1 \mem_reg_93][5  ( .D(D_5), .E(n6251), .C(wclk), .QN(n3907) );
  DFE1 \mem_reg_93][4  ( .D(D_4), .E(n6251), .C(wclk), .QN(n3908) );
  DFE1 \mem_reg_93][3  ( .D(D_3), .E(n6251), .C(wclk), .QN(n3909) );
  DFE1 \mem_reg_93][2  ( .D(D_2), .E(n6251), .C(wclk), .QN(n3910) );
  DFE1 \mem_reg_93][1  ( .D(D_1), .E(n6251), .C(wclk), .QN(n3911) );
  DFE1 \mem_reg_93][0  ( .D(D_0), .E(n6251), .C(wclk), .QN(n3912) );
  DFE1 \mem_reg_92][23  ( .D(D_23), .E(n6250), .C(wclk), .QN(n3913) );
  DFE1 \mem_reg_92][22  ( .D(D_22), .E(n6250), .C(wclk), .QN(n3914) );
  DFE1 \mem_reg_92][21  ( .D(D_21), .E(n6250), .C(wclk), .QN(n3915) );
  DFE1 \mem_reg_92][20  ( .D(D_20), .E(n6250), .C(wclk), .QN(n3916) );
  DFE1 \mem_reg_92][19  ( .D(D_19), .E(n6250), .C(wclk), .QN(n3917) );
  DFE1 \mem_reg_92][18  ( .D(D_18), .E(n6250), .C(wclk), .QN(n3918) );
  DFE1 \mem_reg_92][17  ( .D(D_17), .E(n6250), .C(wclk), .QN(n3919) );
  DFE1 \mem_reg_92][16  ( .D(D_16), .E(n6250), .C(wclk), .QN(n3920) );
  DFE1 \mem_reg_92][15  ( .D(D_15), .E(n6250), .C(wclk), .QN(n3921) );
  DFE1 \mem_reg_92][14  ( .D(D_14), .E(n6250), .C(wclk), .QN(n3922) );
  DFE1 \mem_reg_92][13  ( .D(D_13), .E(n6250), .C(wclk), .QN(n3923) );
  DFE1 \mem_reg_92][12  ( .D(D_12), .E(n6250), .C(wclk), .QN(n3924) );
  DFE1 \mem_reg_92][11  ( .D(D_11), .E(n6250), .C(wclk), .QN(n3925) );
  DFE1 \mem_reg_92][10  ( .D(D_10), .E(n6250), .C(wclk), .QN(n3926) );
  DFE1 \mem_reg_92][9  ( .D(D_9), .E(n6250), .C(wclk), .QN(n3927) );
  DFE1 \mem_reg_92][8  ( .D(D_8), .E(n6250), .C(wclk), .QN(n3928) );
  DFE1 \mem_reg_92][7  ( .D(D_7), .E(n6250), .C(wclk), .QN(n3929) );
  DFE1 \mem_reg_92][6  ( .D(D_6), .E(n6250), .C(wclk), .QN(n3930) );
  DFE1 \mem_reg_92][5  ( .D(D_5), .E(n6250), .C(wclk), .QN(n3931) );
  DFE1 \mem_reg_92][4  ( .D(D_4), .E(n6250), .C(wclk), .QN(n3932) );
  DFE1 \mem_reg_92][3  ( .D(D_3), .E(n6250), .C(wclk), .QN(n3933) );
  DFE1 \mem_reg_92][2  ( .D(D_2), .E(n6250), .C(wclk), .QN(n3934) );
  DFE1 \mem_reg_92][1  ( .D(D_1), .E(n6250), .C(wclk), .QN(n3935) );
  DFE1 \mem_reg_92][0  ( .D(D_0), .E(n6250), .C(wclk), .QN(n3936) );
  DFE1 \mem_reg_91][23  ( .D(D_23), .E(n6249), .C(wclk), .QN(n3937) );
  DFE1 \mem_reg_91][22  ( .D(D_22), .E(n6249), .C(wclk), .QN(n3938) );
  DFE1 \mem_reg_91][21  ( .D(D_21), .E(n6249), .C(wclk), .QN(n3939) );
  DFE1 \mem_reg_91][20  ( .D(D_20), .E(n6249), .C(wclk), .QN(n3940) );
  DFE1 \mem_reg_91][19  ( .D(D_19), .E(n6249), .C(wclk), .QN(n3941) );
  DFE1 \mem_reg_91][18  ( .D(D_18), .E(n6249), .C(wclk), .QN(n3942) );
  DFE1 \mem_reg_91][17  ( .D(D_17), .E(n6249), .C(wclk), .QN(n3943) );
  DFE1 \mem_reg_91][16  ( .D(D_16), .E(n6249), .C(wclk), .QN(n3944) );
  DFE1 \mem_reg_91][15  ( .D(D_15), .E(n6249), .C(wclk), .QN(n3945) );
  DFE1 \mem_reg_91][14  ( .D(D_14), .E(n6249), .C(wclk), .QN(n3946) );
  DFE1 \mem_reg_91][13  ( .D(D_13), .E(n6249), .C(wclk), .QN(n3947) );
  DFE1 \mem_reg_91][12  ( .D(D_12), .E(n6249), .C(wclk), .QN(n3948) );
  DFE1 \mem_reg_91][11  ( .D(D_11), .E(n6249), .C(wclk), .QN(n3949) );
  DFE1 \mem_reg_91][10  ( .D(D_10), .E(n6249), .C(wclk), .QN(n3950) );
  DFE1 \mem_reg_91][9  ( .D(D_9), .E(n6249), .C(wclk), .QN(n3951) );
  DFE1 \mem_reg_91][8  ( .D(D_8), .E(n6249), .C(wclk), .QN(n3952) );
  DFE1 \mem_reg_91][7  ( .D(D_7), .E(n6249), .C(wclk), .QN(n3953) );
  DFE1 \mem_reg_91][6  ( .D(D_6), .E(n6249), .C(wclk), .QN(n3954) );
  DFE1 \mem_reg_91][5  ( .D(D_5), .E(n6249), .C(wclk), .QN(n3955) );
  DFE1 \mem_reg_91][4  ( .D(D_4), .E(n6249), .C(wclk), .QN(n3956) );
  DFE1 \mem_reg_91][3  ( .D(D_3), .E(n6249), .C(wclk), .QN(n3957) );
  DFE1 \mem_reg_91][2  ( .D(D_2), .E(n6249), .C(wclk), .QN(n3958) );
  DFE1 \mem_reg_91][1  ( .D(D_1), .E(n6249), .C(wclk), .QN(n3959) );
  DFE1 \mem_reg_91][0  ( .D(D_0), .E(n6249), .C(wclk), .QN(n3960) );
  DFE1 \mem_reg_90][23  ( .D(D_23), .E(n6248), .C(wclk), .QN(n3961) );
  DFE1 \mem_reg_90][22  ( .D(D_22), .E(n6248), .C(wclk), .QN(n3962) );
  DFE1 \mem_reg_90][21  ( .D(D_21), .E(n6248), .C(wclk), .QN(n3963) );
  DFE1 \mem_reg_90][20  ( .D(D_20), .E(n6248), .C(wclk), .QN(n3964) );
  DFE1 \mem_reg_90][19  ( .D(D_19), .E(n6248), .C(wclk), .QN(n3965) );
  DFE1 \mem_reg_90][18  ( .D(D_18), .E(n6248), .C(wclk), .QN(n3966) );
  DFE1 \mem_reg_90][17  ( .D(D_17), .E(n6248), .C(wclk), .QN(n3967) );
  DFE1 \mem_reg_90][16  ( .D(D_16), .E(n6248), .C(wclk), .QN(n3968) );
  DFE1 \mem_reg_90][15  ( .D(D_15), .E(n6248), .C(wclk), .QN(n3969) );
  DFE1 \mem_reg_90][14  ( .D(D_14), .E(n6248), .C(wclk), .QN(n3970) );
  DFE1 \mem_reg_90][13  ( .D(D_13), .E(n6248), .C(wclk), .QN(n3971) );
  DFE1 \mem_reg_90][12  ( .D(D_12), .E(n6248), .C(wclk), .QN(n3972) );
  DFE1 \mem_reg_90][11  ( .D(D_11), .E(n6248), .C(wclk), .QN(n3973) );
  DFE1 \mem_reg_90][10  ( .D(D_10), .E(n6248), .C(wclk), .QN(n3974) );
  DFE1 \mem_reg_90][9  ( .D(D_9), .E(n6248), .C(wclk), .QN(n3975) );
  DFE1 \mem_reg_90][8  ( .D(D_8), .E(n6248), .C(wclk), .QN(n3976) );
  DFE1 \mem_reg_90][7  ( .D(D_7), .E(n6248), .C(wclk), .QN(n3977) );
  DFE1 \mem_reg_90][6  ( .D(D_6), .E(n6248), .C(wclk), .QN(n3978) );
  DFE1 \mem_reg_90][5  ( .D(D_5), .E(n6248), .C(wclk), .QN(n3979) );
  DFE1 \mem_reg_90][4  ( .D(D_4), .E(n6248), .C(wclk), .QN(n3980) );
  DFE1 \mem_reg_90][3  ( .D(D_3), .E(n6248), .C(wclk), .QN(n3981) );
  DFE1 \mem_reg_90][2  ( .D(D_2), .E(n6248), .C(wclk), .QN(n3982) );
  DFE1 \mem_reg_90][1  ( .D(D_1), .E(n6248), .C(wclk), .QN(n3983) );
  DFE1 \mem_reg_90][0  ( .D(D_0), .E(n6248), .C(wclk), .QN(n3984) );
  DFE1 \mem_reg_89][23  ( .D(D_23), .E(n6247), .C(wclk), .QN(n3985) );
  DFE1 \mem_reg_89][22  ( .D(D_22), .E(n6247), .C(wclk), .QN(n3986) );
  DFE1 \mem_reg_89][21  ( .D(D_21), .E(n6247), .C(wclk), .QN(n3987) );
  DFE1 \mem_reg_89][20  ( .D(D_20), .E(n6247), .C(wclk), .QN(n3988) );
  DFE1 \mem_reg_89][19  ( .D(D_19), .E(n6247), .C(wclk), .QN(n3989) );
  DFE1 \mem_reg_89][18  ( .D(D_18), .E(n6247), .C(wclk), .QN(n3990) );
  DFE1 \mem_reg_89][17  ( .D(D_17), .E(n6247), .C(wclk), .QN(n3991) );
  DFE1 \mem_reg_89][16  ( .D(D_16), .E(n6247), .C(wclk), .QN(n3992) );
  DFE1 \mem_reg_89][15  ( .D(D_15), .E(n6247), .C(wclk), .QN(n3993) );
  DFE1 \mem_reg_89][14  ( .D(D_14), .E(n6247), .C(wclk), .QN(n3994) );
  DFE1 \mem_reg_89][13  ( .D(D_13), .E(n6247), .C(wclk), .QN(n3995) );
  DFE1 \mem_reg_89][12  ( .D(D_12), .E(n6247), .C(wclk), .QN(n3996) );
  DFE1 \mem_reg_89][11  ( .D(D_11), .E(n6247), .C(wclk), .QN(n3997) );
  DFE1 \mem_reg_89][10  ( .D(D_10), .E(n6247), .C(wclk), .QN(n3998) );
  DFE1 \mem_reg_89][9  ( .D(D_9), .E(n6247), .C(wclk), .QN(n3999) );
  DFE1 \mem_reg_89][8  ( .D(D_8), .E(n6247), .C(wclk), .QN(n4000) );
  DFE1 \mem_reg_89][7  ( .D(D_7), .E(n6247), .C(wclk), .QN(n4001) );
  DFE1 \mem_reg_89][6  ( .D(D_6), .E(n6247), .C(wclk), .QN(n4002) );
  DFE1 \mem_reg_89][5  ( .D(D_5), .E(n6247), .C(wclk), .QN(n4003) );
  DFE1 \mem_reg_89][4  ( .D(D_4), .E(n6247), .C(wclk), .QN(n4004) );
  DFE1 \mem_reg_89][3  ( .D(D_3), .E(n6247), .C(wclk), .QN(n4005) );
  DFE1 \mem_reg_89][2  ( .D(D_2), .E(n6247), .C(wclk), .QN(n4006) );
  DFE1 \mem_reg_89][1  ( .D(D_1), .E(n6247), .C(wclk), .QN(n4007) );
  DFE1 \mem_reg_89][0  ( .D(D_0), .E(n6247), .C(wclk), .QN(n4008) );
  DFE1 \mem_reg_88][23  ( .D(D_23), .E(n6246), .C(wclk), .QN(n4009) );
  DFE1 \mem_reg_88][22  ( .D(D_22), .E(n6246), .C(wclk), .QN(n4010) );
  DFE1 \mem_reg_88][21  ( .D(D_21), .E(n6246), .C(wclk), .QN(n4011) );
  DFE1 \mem_reg_88][20  ( .D(D_20), .E(n6246), .C(wclk), .QN(n4012) );
  DFE1 \mem_reg_88][19  ( .D(D_19), .E(n6246), .C(wclk), .QN(n4013) );
  DFE1 \mem_reg_88][18  ( .D(D_18), .E(n6246), .C(wclk), .QN(n4014) );
  DFE1 \mem_reg_88][17  ( .D(D_17), .E(n6246), .C(wclk), .QN(n4015) );
  DFE1 \mem_reg_88][16  ( .D(D_16), .E(n6246), .C(wclk), .QN(n4016) );
  DFE1 \mem_reg_88][15  ( .D(D_15), .E(n6246), .C(wclk), .QN(n4017) );
  DFE1 \mem_reg_88][14  ( .D(D_14), .E(n6246), .C(wclk), .QN(n4018) );
  DFE1 \mem_reg_88][13  ( .D(D_13), .E(n6246), .C(wclk), .QN(n4019) );
  DFE1 \mem_reg_88][12  ( .D(D_12), .E(n6246), .C(wclk), .QN(n4020) );
  DFE1 \mem_reg_88][11  ( .D(D_11), .E(n6246), .C(wclk), .QN(n4021) );
  DFE1 \mem_reg_88][10  ( .D(D_10), .E(n6246), .C(wclk), .QN(n4022) );
  DFE1 \mem_reg_88][9  ( .D(D_9), .E(n6246), .C(wclk), .QN(n4023) );
  DFE1 \mem_reg_88][8  ( .D(D_8), .E(n6246), .C(wclk), .QN(n4024) );
  DFE1 \mem_reg_88][7  ( .D(D_7), .E(n6246), .C(wclk), .QN(n4025) );
  DFE1 \mem_reg_88][6  ( .D(D_6), .E(n6246), .C(wclk), .QN(n4026) );
  DFE1 \mem_reg_88][5  ( .D(D_5), .E(n6246), .C(wclk), .QN(n4027) );
  DFE1 \mem_reg_88][4  ( .D(D_4), .E(n6246), .C(wclk), .QN(n4028) );
  DFE1 \mem_reg_88][3  ( .D(D_3), .E(n6246), .C(wclk), .QN(n4029) );
  DFE1 \mem_reg_88][2  ( .D(D_2), .E(n6246), .C(wclk), .QN(n4030) );
  DFE1 \mem_reg_88][1  ( .D(D_1), .E(n6246), .C(wclk), .QN(n4031) );
  DFE1 \mem_reg_88][0  ( .D(D_0), .E(n6246), .C(wclk), .QN(n4032) );
  DFE1 \mem_reg_87][23  ( .D(D_23), .E(n6245), .C(wclk), .QN(n4033) );
  DFE1 \mem_reg_87][22  ( .D(D_22), .E(n6245), .C(wclk), .QN(n4034) );
  DFE1 \mem_reg_87][21  ( .D(D_21), .E(n6245), .C(wclk), .QN(n4035) );
  DFE1 \mem_reg_87][20  ( .D(D_20), .E(n6245), .C(wclk), .QN(n4036) );
  DFE1 \mem_reg_87][19  ( .D(D_19), .E(n6245), .C(wclk), .QN(n4037) );
  DFE1 \mem_reg_87][18  ( .D(D_18), .E(n6245), .C(wclk), .QN(n4038) );
  DFE1 \mem_reg_87][17  ( .D(D_17), .E(n6245), .C(wclk), .QN(n4039) );
  DFE1 \mem_reg_87][16  ( .D(D_16), .E(n6245), .C(wclk), .QN(n4040) );
  DFE1 \mem_reg_87][15  ( .D(D_15), .E(n6245), .C(wclk), .QN(n4041) );
  DFE1 \mem_reg_87][14  ( .D(D_14), .E(n6245), .C(wclk), .QN(n4042) );
  DFE1 \mem_reg_87][13  ( .D(D_13), .E(n6245), .C(wclk), .QN(n4043) );
  DFE1 \mem_reg_87][12  ( .D(D_12), .E(n6245), .C(wclk), .QN(n4044) );
  DFE1 \mem_reg_87][11  ( .D(D_11), .E(n6245), .C(wclk), .QN(n4045) );
  DFE1 \mem_reg_87][10  ( .D(D_10), .E(n6245), .C(wclk), .QN(n4046) );
  DFE1 \mem_reg_87][9  ( .D(D_9), .E(n6245), .C(wclk), .QN(n4047) );
  DFE1 \mem_reg_87][8  ( .D(D_8), .E(n6245), .C(wclk), .QN(n4048) );
  DFE1 \mem_reg_87][7  ( .D(D_7), .E(n6245), .C(wclk), .QN(n4049) );
  DFE1 \mem_reg_87][6  ( .D(D_6), .E(n6245), .C(wclk), .QN(n4050) );
  DFE1 \mem_reg_87][5  ( .D(D_5), .E(n6245), .C(wclk), .QN(n4051) );
  DFE1 \mem_reg_87][4  ( .D(D_4), .E(n6245), .C(wclk), .QN(n4052) );
  DFE1 \mem_reg_87][3  ( .D(D_3), .E(n6245), .C(wclk), .QN(n4053) );
  DFE1 \mem_reg_87][2  ( .D(D_2), .E(n6245), .C(wclk), .QN(n4054) );
  DFE1 \mem_reg_87][1  ( .D(D_1), .E(n6245), .C(wclk), .QN(n4055) );
  DFE1 \mem_reg_87][0  ( .D(D_0), .E(n6245), .C(wclk), .QN(n4056) );
  DFE1 \mem_reg_86][23  ( .D(D_23), .E(n6244), .C(wclk), .QN(n4057) );
  DFE1 \mem_reg_86][22  ( .D(D_22), .E(n6244), .C(wclk), .QN(n4058) );
  DFE1 \mem_reg_86][21  ( .D(D_21), .E(n6244), .C(wclk), .QN(n4059) );
  DFE1 \mem_reg_86][20  ( .D(D_20), .E(n6244), .C(wclk), .QN(n4060) );
  DFE1 \mem_reg_86][19  ( .D(D_19), .E(n6244), .C(wclk), .QN(n4061) );
  DFE1 \mem_reg_86][18  ( .D(D_18), .E(n6244), .C(wclk), .QN(n4062) );
  DFE1 \mem_reg_86][17  ( .D(D_17), .E(n6244), .C(wclk), .QN(n4063) );
  DFE1 \mem_reg_86][16  ( .D(D_16), .E(n6244), .C(wclk), .QN(n4064) );
  DFE1 \mem_reg_86][15  ( .D(D_15), .E(n6244), .C(wclk), .QN(n4065) );
  DFE1 \mem_reg_86][14  ( .D(D_14), .E(n6244), .C(wclk), .QN(n4066) );
  DFE1 \mem_reg_86][13  ( .D(D_13), .E(n6244), .C(wclk), .QN(n4067) );
  DFE1 \mem_reg_86][12  ( .D(D_12), .E(n6244), .C(wclk), .QN(n4068) );
  DFE1 \mem_reg_86][11  ( .D(D_11), .E(n6244), .C(wclk), .QN(n4069) );
  DFE1 \mem_reg_86][10  ( .D(D_10), .E(n6244), .C(wclk), .QN(n4070) );
  DFE1 \mem_reg_86][9  ( .D(D_9), .E(n6244), .C(wclk), .QN(n4071) );
  DFE1 \mem_reg_86][8  ( .D(D_8), .E(n6244), .C(wclk), .QN(n4072) );
  DFE1 \mem_reg_86][7  ( .D(D_7), .E(n6244), .C(wclk), .QN(n4073) );
  DFE1 \mem_reg_86][6  ( .D(D_6), .E(n6244), .C(wclk), .QN(n4074) );
  DFE1 \mem_reg_86][5  ( .D(D_5), .E(n6244), .C(wclk), .QN(n4075) );
  DFE1 \mem_reg_86][4  ( .D(D_4), .E(n6244), .C(wclk), .QN(n4076) );
  DFE1 \mem_reg_86][3  ( .D(D_3), .E(n6244), .C(wclk), .QN(n4077) );
  DFE1 \mem_reg_86][2  ( .D(D_2), .E(n6244), .C(wclk), .QN(n4078) );
  DFE1 \mem_reg_86][1  ( .D(D_1), .E(n6244), .C(wclk), .QN(n4079) );
  DFE1 \mem_reg_86][0  ( .D(D_0), .E(n6244), .C(wclk), .QN(n4080) );
  DFE1 \mem_reg_85][23  ( .D(D_23), .E(n6243), .C(wclk), .QN(n4081) );
  DFE1 \mem_reg_85][22  ( .D(D_22), .E(n6243), .C(wclk), .QN(n4082) );
  DFE1 \mem_reg_85][21  ( .D(D_21), .E(n6243), .C(wclk), .QN(n4083) );
  DFE1 \mem_reg_85][20  ( .D(D_20), .E(n6243), .C(wclk), .QN(n4084) );
  DFE1 \mem_reg_85][19  ( .D(D_19), .E(n6243), .C(wclk), .QN(n4085) );
  DFE1 \mem_reg_85][18  ( .D(D_18), .E(n6243), .C(wclk), .QN(n4086) );
  DFE1 \mem_reg_85][17  ( .D(D_17), .E(n6243), .C(wclk), .QN(n4087) );
  DFE1 \mem_reg_85][16  ( .D(D_16), .E(n6243), .C(wclk), .QN(n4088) );
  DFE1 \mem_reg_85][15  ( .D(D_15), .E(n6243), .C(wclk), .QN(n4089) );
  DFE1 \mem_reg_85][14  ( .D(D_14), .E(n6243), .C(wclk), .QN(n4090) );
  DFE1 \mem_reg_85][13  ( .D(D_13), .E(n6243), .C(wclk), .QN(n4091) );
  DFE1 \mem_reg_85][12  ( .D(D_12), .E(n6243), .C(wclk), .QN(n4092) );
  DFE1 \mem_reg_85][11  ( .D(D_11), .E(n6243), .C(wclk), .QN(n4093) );
  DFE1 \mem_reg_85][10  ( .D(D_10), .E(n6243), .C(wclk), .QN(n4094) );
  DFE1 \mem_reg_85][9  ( .D(D_9), .E(n6243), .C(wclk), .QN(n4095) );
  DFE1 \mem_reg_85][8  ( .D(D_8), .E(n6243), .C(wclk), .QN(n4096) );
  DFE1 \mem_reg_85][7  ( .D(D_7), .E(n6243), .C(wclk), .QN(n4097) );
  DFE1 \mem_reg_85][6  ( .D(D_6), .E(n6243), .C(wclk), .QN(n4098) );
  DFE1 \mem_reg_85][5  ( .D(D_5), .E(n6243), .C(wclk), .QN(n4099) );
  DFE1 \mem_reg_85][4  ( .D(D_4), .E(n6243), .C(wclk), .QN(n4100) );
  DFE1 \mem_reg_85][3  ( .D(D_3), .E(n6243), .C(wclk), .QN(n4101) );
  DFE1 \mem_reg_85][2  ( .D(D_2), .E(n6243), .C(wclk), .QN(n4102) );
  DFE1 \mem_reg_85][1  ( .D(D_1), .E(n6243), .C(wclk), .QN(n4103) );
  DFE1 \mem_reg_85][0  ( .D(D_0), .E(n6243), .C(wclk), .QN(n4104) );
  DFE1 \mem_reg_84][23  ( .D(D_23), .E(n6242), .C(wclk), .QN(n4105) );
  DFE1 \mem_reg_84][22  ( .D(D_22), .E(n6242), .C(wclk), .QN(n4106) );
  DFE1 \mem_reg_84][21  ( .D(D_21), .E(n6242), .C(wclk), .QN(n4107) );
  DFE1 \mem_reg_84][20  ( .D(D_20), .E(n6242), .C(wclk), .QN(n4108) );
  DFE1 \mem_reg_84][19  ( .D(D_19), .E(n6242), .C(wclk), .QN(n4109) );
  DFE1 \mem_reg_84][18  ( .D(D_18), .E(n6242), .C(wclk), .QN(n4110) );
  DFE1 \mem_reg_84][17  ( .D(D_17), .E(n6242), .C(wclk), .QN(n4111) );
  DFE1 \mem_reg_84][16  ( .D(D_16), .E(n6242), .C(wclk), .QN(n4112) );
  DFE1 \mem_reg_84][15  ( .D(D_15), .E(n6242), .C(wclk), .QN(n4113) );
  DFE1 \mem_reg_84][14  ( .D(D_14), .E(n6242), .C(wclk), .QN(n4114) );
  DFE1 \mem_reg_84][13  ( .D(D_13), .E(n6242), .C(wclk), .QN(n4115) );
  DFE1 \mem_reg_84][12  ( .D(D_12), .E(n6242), .C(wclk), .QN(n4116) );
  DFE1 \mem_reg_84][11  ( .D(D_11), .E(n6242), .C(wclk), .QN(n4117) );
  DFE1 \mem_reg_84][10  ( .D(D_10), .E(n6242), .C(wclk), .QN(n4118) );
  DFE1 \mem_reg_84][9  ( .D(D_9), .E(n6242), .C(wclk), .QN(n4119) );
  DFE1 \mem_reg_84][8  ( .D(D_8), .E(n6242), .C(wclk), .QN(n4120) );
  DFE1 \mem_reg_84][7  ( .D(D_7), .E(n6242), .C(wclk), .QN(n4121) );
  DFE1 \mem_reg_84][6  ( .D(D_6), .E(n6242), .C(wclk), .QN(n4122) );
  DFE1 \mem_reg_84][5  ( .D(D_5), .E(n6242), .C(wclk), .QN(n4123) );
  DFE1 \mem_reg_84][4  ( .D(D_4), .E(n6242), .C(wclk), .QN(n4124) );
  DFE1 \mem_reg_84][3  ( .D(D_3), .E(n6242), .C(wclk), .QN(n4125) );
  DFE1 \mem_reg_84][2  ( .D(D_2), .E(n6242), .C(wclk), .QN(n4126) );
  DFE1 \mem_reg_84][1  ( .D(D_1), .E(n6242), .C(wclk), .QN(n4127) );
  DFE1 \mem_reg_84][0  ( .D(D_0), .E(n6242), .C(wclk), .QN(n4128) );
  DFE1 \mem_reg_83][23  ( .D(D_23), .E(n6240), .C(wclk), .QN(n4129) );
  DFE1 \mem_reg_83][22  ( .D(D_22), .E(n6240), .C(wclk), .QN(n4130) );
  DFE1 \mem_reg_83][21  ( .D(D_21), .E(n6240), .C(wclk), .QN(n4131) );
  DFE1 \mem_reg_83][20  ( .D(D_20), .E(n6240), .C(wclk), .QN(n4132) );
  DFE1 \mem_reg_83][19  ( .D(D_19), .E(n6240), .C(wclk), .QN(n4133) );
  DFE1 \mem_reg_83][18  ( .D(D_18), .E(n6240), .C(wclk), .QN(n4134) );
  DFE1 \mem_reg_83][17  ( .D(D_17), .E(n6240), .C(wclk), .QN(n4135) );
  DFE1 \mem_reg_83][16  ( .D(D_16), .E(n6240), .C(wclk), .QN(n4136) );
  DFE1 \mem_reg_83][15  ( .D(D_15), .E(n6240), .C(wclk), .QN(n4137) );
  DFE1 \mem_reg_83][14  ( .D(D_14), .E(n6240), .C(wclk), .QN(n4138) );
  DFE1 \mem_reg_83][13  ( .D(D_13), .E(n6240), .C(wclk), .QN(n4139) );
  DFE1 \mem_reg_83][12  ( .D(D_12), .E(n6240), .C(wclk), .QN(n4140) );
  DFE1 \mem_reg_83][11  ( .D(D_11), .E(n6240), .C(wclk), .QN(n4141) );
  DFE1 \mem_reg_83][10  ( .D(D_10), .E(n6240), .C(wclk), .QN(n4142) );
  DFE1 \mem_reg_83][9  ( .D(D_9), .E(n6240), .C(wclk), .QN(n4143) );
  DFE1 \mem_reg_83][8  ( .D(D_8), .E(n6240), .C(wclk), .QN(n4144) );
  DFE1 \mem_reg_83][7  ( .D(D_7), .E(n6240), .C(wclk), .QN(n4145) );
  DFE1 \mem_reg_83][6  ( .D(D_6), .E(n6240), .C(wclk), .QN(n4146) );
  DFE1 \mem_reg_83][5  ( .D(D_5), .E(n6240), .C(wclk), .QN(n4147) );
  DFE1 \mem_reg_83][4  ( .D(D_4), .E(n6240), .C(wclk), .QN(n4148) );
  DFE1 \mem_reg_83][3  ( .D(D_3), .E(n6240), .C(wclk), .QN(n4149) );
  DFE1 \mem_reg_83][2  ( .D(D_2), .E(n6240), .C(wclk), .QN(n4150) );
  DFE1 \mem_reg_83][1  ( .D(D_1), .E(n6240), .C(wclk), .QN(n4151) );
  DFE1 \mem_reg_83][0  ( .D(D_0), .E(n6240), .C(wclk), .QN(n4152) );
  DFE1 \mem_reg_82][23  ( .D(D_23), .E(n6239), .C(wclk), .QN(n4153) );
  DFE1 \mem_reg_82][22  ( .D(D_22), .E(n6239), .C(wclk), .QN(n4154) );
  DFE1 \mem_reg_82][21  ( .D(D_21), .E(n6239), .C(wclk), .QN(n4155) );
  DFE1 \mem_reg_82][20  ( .D(D_20), .E(n6239), .C(wclk), .QN(n4156) );
  DFE1 \mem_reg_82][19  ( .D(D_19), .E(n6239), .C(wclk), .QN(n4157) );
  DFE1 \mem_reg_82][18  ( .D(D_18), .E(n6239), .C(wclk), .QN(n4158) );
  DFE1 \mem_reg_82][17  ( .D(D_17), .E(n6239), .C(wclk), .QN(n4159) );
  DFE1 \mem_reg_82][16  ( .D(D_16), .E(n6239), .C(wclk), .QN(n4160) );
  DFE1 \mem_reg_82][15  ( .D(D_15), .E(n6239), .C(wclk), .QN(n4161) );
  DFE1 \mem_reg_82][14  ( .D(D_14), .E(n6239), .C(wclk), .QN(n4162) );
  DFE1 \mem_reg_82][13  ( .D(D_13), .E(n6239), .C(wclk), .QN(n4163) );
  DFE1 \mem_reg_82][12  ( .D(D_12), .E(n6239), .C(wclk), .QN(n4164) );
  DFE1 \mem_reg_82][11  ( .D(D_11), .E(n6239), .C(wclk), .QN(n4165) );
  DFE1 \mem_reg_82][10  ( .D(D_10), .E(n6239), .C(wclk), .QN(n4166) );
  DFE1 \mem_reg_82][9  ( .D(D_9), .E(n6239), .C(wclk), .QN(n4167) );
  DFE1 \mem_reg_82][8  ( .D(D_8), .E(n6239), .C(wclk), .QN(n4168) );
  DFE1 \mem_reg_82][7  ( .D(D_7), .E(n6239), .C(wclk), .QN(n4169) );
  DFE1 \mem_reg_82][6  ( .D(D_6), .E(n6239), .C(wclk), .QN(n4170) );
  DFE1 \mem_reg_82][5  ( .D(D_5), .E(n6239), .C(wclk), .QN(n4171) );
  DFE1 \mem_reg_82][4  ( .D(D_4), .E(n6239), .C(wclk), .QN(n4172) );
  DFE1 \mem_reg_82][3  ( .D(D_3), .E(n6239), .C(wclk), .QN(n4173) );
  DFE1 \mem_reg_82][2  ( .D(D_2), .E(n6239), .C(wclk), .QN(n4174) );
  DFE1 \mem_reg_82][1  ( .D(D_1), .E(n6239), .C(wclk), .QN(n4175) );
  DFE1 \mem_reg_82][0  ( .D(D_0), .E(n6239), .C(wclk), .QN(n4176) );
  DFE1 \mem_reg_81][23  ( .D(D_23), .E(n6238), .C(wclk), .QN(n4177) );
  DFE1 \mem_reg_81][22  ( .D(D_22), .E(n6238), .C(wclk), .QN(n4178) );
  DFE1 \mem_reg_81][21  ( .D(D_21), .E(n6238), .C(wclk), .QN(n4179) );
  DFE1 \mem_reg_81][20  ( .D(D_20), .E(n6238), .C(wclk), .QN(n4180) );
  DFE1 \mem_reg_81][19  ( .D(D_19), .E(n6238), .C(wclk), .QN(n4181) );
  DFE1 \mem_reg_81][18  ( .D(D_18), .E(n6238), .C(wclk), .QN(n4182) );
  DFE1 \mem_reg_81][17  ( .D(D_17), .E(n6238), .C(wclk), .QN(n4183) );
  DFE1 \mem_reg_81][16  ( .D(D_16), .E(n6238), .C(wclk), .QN(n4184) );
  DFE1 \mem_reg_81][15  ( .D(D_15), .E(n6238), .C(wclk), .QN(n4185) );
  DFE1 \mem_reg_81][14  ( .D(D_14), .E(n6238), .C(wclk), .QN(n4186) );
  DFE1 \mem_reg_81][13  ( .D(D_13), .E(n6238), .C(wclk), .QN(n4187) );
  DFE1 \mem_reg_81][12  ( .D(D_12), .E(n6238), .C(wclk), .QN(n4188) );
  DFE1 \mem_reg_81][11  ( .D(D_11), .E(n6238), .C(wclk), .QN(n4189) );
  DFE1 \mem_reg_81][10  ( .D(D_10), .E(n6238), .C(wclk), .QN(n4190) );
  DFE1 \mem_reg_81][9  ( .D(D_9), .E(n6238), .C(wclk), .QN(n4191) );
  DFE1 \mem_reg_81][8  ( .D(D_8), .E(n6238), .C(wclk), .QN(n4192) );
  DFE1 \mem_reg_81][7  ( .D(D_7), .E(n6238), .C(wclk), .QN(n4193) );
  DFE1 \mem_reg_81][6  ( .D(D_6), .E(n6238), .C(wclk), .QN(n4194) );
  DFE1 \mem_reg_81][5  ( .D(D_5), .E(n6238), .C(wclk), .QN(n4195) );
  DFE1 \mem_reg_81][4  ( .D(D_4), .E(n6238), .C(wclk), .QN(n4196) );
  DFE1 \mem_reg_81][3  ( .D(D_3), .E(n6238), .C(wclk), .QN(n4197) );
  DFE1 \mem_reg_81][2  ( .D(D_2), .E(n6238), .C(wclk), .QN(n4198) );
  DFE1 \mem_reg_81][1  ( .D(D_1), .E(n6238), .C(wclk), .QN(n4199) );
  DFE1 \mem_reg_81][0  ( .D(D_0), .E(n6238), .C(wclk), .QN(n4200) );
  DFE1 \mem_reg_80][23  ( .D(D_23), .E(n6236), .C(wclk), .QN(n4201) );
  DFE1 \mem_reg_80][22  ( .D(D_22), .E(n6236), .C(wclk), .QN(n4202) );
  DFE1 \mem_reg_80][21  ( .D(D_21), .E(n6236), .C(wclk), .QN(n4203) );
  DFE1 \mem_reg_80][20  ( .D(D_20), .E(n6236), .C(wclk), .QN(n4204) );
  DFE1 \mem_reg_80][19  ( .D(D_19), .E(n6236), .C(wclk), .QN(n4205) );
  DFE1 \mem_reg_80][18  ( .D(D_18), .E(n6236), .C(wclk), .QN(n4206) );
  DFE1 \mem_reg_80][17  ( .D(D_17), .E(n6236), .C(wclk), .QN(n4207) );
  DFE1 \mem_reg_80][16  ( .D(D_16), .E(n6236), .C(wclk), .QN(n4208) );
  DFE1 \mem_reg_80][15  ( .D(D_15), .E(n6236), .C(wclk), .QN(n4209) );
  DFE1 \mem_reg_80][14  ( .D(D_14), .E(n6236), .C(wclk), .QN(n4210) );
  DFE1 \mem_reg_80][13  ( .D(D_13), .E(n6236), .C(wclk), .QN(n4211) );
  DFE1 \mem_reg_80][12  ( .D(D_12), .E(n6236), .C(wclk), .QN(n4212) );
  DFE1 \mem_reg_80][11  ( .D(D_11), .E(n6236), .C(wclk), .QN(n4213) );
  DFE1 \mem_reg_80][10  ( .D(D_10), .E(n6236), .C(wclk), .QN(n4214) );
  DFE1 \mem_reg_80][9  ( .D(D_9), .E(n6236), .C(wclk), .QN(n4215) );
  DFE1 \mem_reg_80][8  ( .D(D_8), .E(n6236), .C(wclk), .QN(n4216) );
  DFE1 \mem_reg_80][7  ( .D(D_7), .E(n6236), .C(wclk), .QN(n4217) );
  DFE1 \mem_reg_80][6  ( .D(D_6), .E(n6236), .C(wclk), .QN(n4218) );
  DFE1 \mem_reg_80][5  ( .D(D_5), .E(n6236), .C(wclk), .QN(n4219) );
  DFE1 \mem_reg_80][4  ( .D(D_4), .E(n6236), .C(wclk), .QN(n4220) );
  DFE1 \mem_reg_80][3  ( .D(D_3), .E(n6236), .C(wclk), .QN(n4221) );
  DFE1 \mem_reg_80][2  ( .D(D_2), .E(n6236), .C(wclk), .QN(n4222) );
  DFE1 \mem_reg_80][1  ( .D(D_1), .E(n6236), .C(wclk), .QN(n4223) );
  DFE1 \mem_reg_80][0  ( .D(D_0), .E(n6236), .C(wclk), .QN(n4224) );
  DFE1 \mem_reg_47][23  ( .D(D_23), .E(n6477), .C(wclk), .QN(n4993) );
  DFE1 \mem_reg_47][22  ( .D(D_22), .E(n6477), .C(wclk), .QN(n4994) );
  DFE1 \mem_reg_47][21  ( .D(D_21), .E(n6477), .C(wclk), .QN(n4995) );
  DFE1 \mem_reg_47][20  ( .D(D_20), .E(n6477), .C(wclk), .QN(n4996) );
  DFE1 \mem_reg_47][19  ( .D(D_19), .E(n6477), .C(wclk), .QN(n4997) );
  DFE1 \mem_reg_47][18  ( .D(D_18), .E(n6477), .C(wclk), .QN(n4998) );
  DFE1 \mem_reg_47][17  ( .D(D_17), .E(n6477), .C(wclk), .QN(n4999) );
  DFE1 \mem_reg_47][16  ( .D(D_16), .E(n6477), .C(wclk), .QN(n5000) );
  DFE1 \mem_reg_47][15  ( .D(D_15), .E(n6477), .C(wclk), .QN(n5001) );
  DFE1 \mem_reg_47][14  ( .D(D_14), .E(n6477), .C(wclk), .QN(n5002) );
  DFE1 \mem_reg_47][13  ( .D(D_13), .E(n6477), .C(wclk), .QN(n5003) );
  DFE1 \mem_reg_47][12  ( .D(D_12), .E(n6477), .C(wclk), .QN(n5004) );
  DFE1 \mem_reg_47][11  ( .D(D_11), .E(n6477), .C(wclk), .QN(n5005) );
  DFE1 \mem_reg_47][10  ( .D(D_10), .E(n6477), .C(wclk), .QN(n5006) );
  DFE1 \mem_reg_47][9  ( .D(D_9), .E(n6477), .C(wclk), .QN(n5007) );
  DFE1 \mem_reg_47][8  ( .D(D_8), .E(n6477), .C(wclk), .QN(n5008) );
  DFE1 \mem_reg_47][7  ( .D(D_7), .E(n6477), .C(wclk), .QN(n5009) );
  DFE1 \mem_reg_47][6  ( .D(D_6), .E(n6477), .C(wclk), .QN(n5010) );
  DFE1 \mem_reg_47][5  ( .D(D_5), .E(n6477), .C(wclk), .QN(n5011) );
  DFE1 \mem_reg_47][4  ( .D(D_4), .E(n6477), .C(wclk), .QN(n5012) );
  DFE1 \mem_reg_47][3  ( .D(D_3), .E(n6477), .C(wclk), .QN(n5013) );
  DFE1 \mem_reg_47][2  ( .D(D_2), .E(n6477), .C(wclk), .QN(n5014) );
  DFE1 \mem_reg_47][1  ( .D(D_1), .E(n6477), .C(wclk), .QN(n5015) );
  DFE1 \mem_reg_47][0  ( .D(D_0), .E(n6477), .C(wclk), .QN(n5016) );
  DFE1 \mem_reg_46][23  ( .D(D_23), .E(n6474), .C(wclk), .QN(n5017) );
  DFE1 \mem_reg_46][22  ( .D(D_22), .E(n6474), .C(wclk), .QN(n5018) );
  DFE1 \mem_reg_46][21  ( .D(D_21), .E(n6474), .C(wclk), .QN(n5019) );
  DFE1 \mem_reg_46][20  ( .D(D_20), .E(n6474), .C(wclk), .QN(n5020) );
  DFE1 \mem_reg_46][19  ( .D(D_19), .E(n6474), .C(wclk), .QN(n5021) );
  DFE1 \mem_reg_46][18  ( .D(D_18), .E(n6474), .C(wclk), .QN(n5022) );
  DFE1 \mem_reg_46][17  ( .D(D_17), .E(n6474), .C(wclk), .QN(n5023) );
  DFE1 \mem_reg_46][16  ( .D(D_16), .E(n6474), .C(wclk), .QN(n5024) );
  DFE1 \mem_reg_46][15  ( .D(D_15), .E(n6474), .C(wclk), .QN(n5025) );
  DFE1 \mem_reg_46][14  ( .D(D_14), .E(n6474), .C(wclk), .QN(n5026) );
  DFE1 \mem_reg_46][13  ( .D(D_13), .E(n6474), .C(wclk), .QN(n5027) );
  DFE1 \mem_reg_46][12  ( .D(D_12), .E(n6474), .C(wclk), .QN(n5028) );
  DFE1 \mem_reg_46][11  ( .D(D_11), .E(n6474), .C(wclk), .QN(n5029) );
  DFE1 \mem_reg_46][10  ( .D(D_10), .E(n6474), .C(wclk), .QN(n5030) );
  DFE1 \mem_reg_46][9  ( .D(D_9), .E(n6474), .C(wclk), .QN(n5031) );
  DFE1 \mem_reg_46][8  ( .D(D_8), .E(n6474), .C(wclk), .QN(n5032) );
  DFE1 \mem_reg_46][7  ( .D(D_7), .E(n6474), .C(wclk), .QN(n5033) );
  DFE1 \mem_reg_46][6  ( .D(D_6), .E(n6474), .C(wclk), .QN(n5034) );
  DFE1 \mem_reg_46][5  ( .D(D_5), .E(n6474), .C(wclk), .QN(n5035) );
  DFE1 \mem_reg_46][4  ( .D(D_4), .E(n6474), .C(wclk), .QN(n5036) );
  DFE1 \mem_reg_46][3  ( .D(D_3), .E(n6474), .C(wclk), .QN(n5037) );
  DFE1 \mem_reg_46][2  ( .D(D_2), .E(n6474), .C(wclk), .QN(n5038) );
  DFE1 \mem_reg_46][1  ( .D(D_1), .E(n6474), .C(wclk), .QN(n5039) );
  DFE1 \mem_reg_46][0  ( .D(D_0), .E(n6474), .C(wclk), .QN(n5040) );
  DFE1 \mem_reg_45][23  ( .D(D_23), .E(n6473), .C(wclk), .QN(n5041) );
  DFE1 \mem_reg_45][22  ( .D(D_22), .E(n6473), .C(wclk), .QN(n5042) );
  DFE1 \mem_reg_45][21  ( .D(D_21), .E(n6473), .C(wclk), .QN(n5043) );
  DFE1 \mem_reg_45][20  ( .D(D_20), .E(n6473), .C(wclk), .QN(n5044) );
  DFE1 \mem_reg_45][19  ( .D(D_19), .E(n6473), .C(wclk), .QN(n5045) );
  DFE1 \mem_reg_45][18  ( .D(D_18), .E(n6473), .C(wclk), .QN(n5046) );
  DFE1 \mem_reg_45][17  ( .D(D_17), .E(n6473), .C(wclk), .QN(n5047) );
  DFE1 \mem_reg_45][16  ( .D(D_16), .E(n6473), .C(wclk), .QN(n5048) );
  DFE1 \mem_reg_45][15  ( .D(D_15), .E(n6473), .C(wclk), .QN(n5049) );
  DFE1 \mem_reg_45][14  ( .D(D_14), .E(n6473), .C(wclk), .QN(n5050) );
  DFE1 \mem_reg_45][13  ( .D(D_13), .E(n6473), .C(wclk), .QN(n5051) );
  DFE1 \mem_reg_45][12  ( .D(D_12), .E(n6473), .C(wclk), .QN(n5052) );
  DFE1 \mem_reg_45][11  ( .D(D_11), .E(n6473), .C(wclk), .QN(n5053) );
  DFE1 \mem_reg_45][10  ( .D(D_10), .E(n6473), .C(wclk), .QN(n5054) );
  DFE1 \mem_reg_45][9  ( .D(D_9), .E(n6473), .C(wclk), .QN(n5055) );
  DFE1 \mem_reg_45][8  ( .D(D_8), .E(n6473), .C(wclk), .QN(n5056) );
  DFE1 \mem_reg_45][7  ( .D(D_7), .E(n6473), .C(wclk), .QN(n5057) );
  DFE1 \mem_reg_45][6  ( .D(D_6), .E(n6473), .C(wclk), .QN(n5058) );
  DFE1 \mem_reg_45][5  ( .D(D_5), .E(n6473), .C(wclk), .QN(n5059) );
  DFE1 \mem_reg_45][4  ( .D(D_4), .E(n6473), .C(wclk), .QN(n5060) );
  DFE1 \mem_reg_45][3  ( .D(D_3), .E(n6473), .C(wclk), .QN(n5061) );
  DFE1 \mem_reg_45][2  ( .D(D_2), .E(n6473), .C(wclk), .QN(n5062) );
  DFE1 \mem_reg_45][1  ( .D(D_1), .E(n6473), .C(wclk), .QN(n5063) );
  DFE1 \mem_reg_45][0  ( .D(D_0), .E(n6473), .C(wclk), .QN(n5064) );
  DFE1 \mem_reg_44][23  ( .D(D_23), .E(n6472), .C(wclk), .QN(n5065) );
  DFE1 \mem_reg_44][22  ( .D(D_22), .E(n6472), .C(wclk), .QN(n5066) );
  DFE1 \mem_reg_44][21  ( .D(D_21), .E(n6472), .C(wclk), .QN(n5067) );
  DFE1 \mem_reg_44][20  ( .D(D_20), .E(n6472), .C(wclk), .QN(n5068) );
  DFE1 \mem_reg_44][19  ( .D(D_19), .E(n6472), .C(wclk), .QN(n5069) );
  DFE1 \mem_reg_44][18  ( .D(D_18), .E(n6472), .C(wclk), .QN(n5070) );
  DFE1 \mem_reg_44][17  ( .D(D_17), .E(n6472), .C(wclk), .QN(n5071) );
  DFE1 \mem_reg_44][16  ( .D(D_16), .E(n6472), .C(wclk), .QN(n5072) );
  DFE1 \mem_reg_44][15  ( .D(D_15), .E(n6472), .C(wclk), .QN(n5073) );
  DFE1 \mem_reg_44][14  ( .D(D_14), .E(n6472), .C(wclk), .QN(n5074) );
  DFE1 \mem_reg_44][13  ( .D(D_13), .E(n6472), .C(wclk), .QN(n5075) );
  DFE1 \mem_reg_44][12  ( .D(D_12), .E(n6472), .C(wclk), .QN(n5076) );
  DFE1 \mem_reg_44][11  ( .D(D_11), .E(n6472), .C(wclk), .QN(n5077) );
  DFE1 \mem_reg_44][10  ( .D(D_10), .E(n6472), .C(wclk), .QN(n5078) );
  DFE1 \mem_reg_44][9  ( .D(D_9), .E(n6472), .C(wclk), .QN(n5079) );
  DFE1 \mem_reg_44][8  ( .D(D_8), .E(n6472), .C(wclk), .QN(n5080) );
  DFE1 \mem_reg_44][7  ( .D(D_7), .E(n6472), .C(wclk), .QN(n5081) );
  DFE1 \mem_reg_44][6  ( .D(D_6), .E(n6472), .C(wclk), .QN(n5082) );
  DFE1 \mem_reg_44][5  ( .D(D_5), .E(n6472), .C(wclk), .QN(n5083) );
  DFE1 \mem_reg_44][4  ( .D(D_4), .E(n6472), .C(wclk), .QN(n5084) );
  DFE1 \mem_reg_44][3  ( .D(D_3), .E(n6472), .C(wclk), .QN(n5085) );
  DFE1 \mem_reg_44][2  ( .D(D_2), .E(n6472), .C(wclk), .QN(n5086) );
  DFE1 \mem_reg_44][1  ( .D(D_1), .E(n6472), .C(wclk), .QN(n5087) );
  DFE1 \mem_reg_44][0  ( .D(D_0), .E(n6472), .C(wclk), .QN(n5088) );
  DFE1 \mem_reg_43][23  ( .D(D_23), .E(n6470), .C(wclk), .QN(n5089) );
  DFE1 \mem_reg_43][22  ( .D(D_22), .E(n6470), .C(wclk), .QN(n5090) );
  DFE1 \mem_reg_43][21  ( .D(D_21), .E(n6470), .C(wclk), .QN(n5091) );
  DFE1 \mem_reg_43][20  ( .D(D_20), .E(n6470), .C(wclk), .QN(n5092) );
  DFE1 \mem_reg_43][19  ( .D(D_19), .E(n6470), .C(wclk), .QN(n5093) );
  DFE1 \mem_reg_43][18  ( .D(D_18), .E(n6470), .C(wclk), .QN(n5094) );
  DFE1 \mem_reg_43][17  ( .D(D_17), .E(n6470), .C(wclk), .QN(n5095) );
  DFE1 \mem_reg_43][16  ( .D(D_16), .E(n6470), .C(wclk), .QN(n5096) );
  DFE1 \mem_reg_43][15  ( .D(D_15), .E(n6470), .C(wclk), .QN(n5097) );
  DFE1 \mem_reg_43][14  ( .D(D_14), .E(n6470), .C(wclk), .QN(n5098) );
  DFE1 \mem_reg_43][13  ( .D(D_13), .E(n6470), .C(wclk), .QN(n5099) );
  DFE1 \mem_reg_43][12  ( .D(D_12), .E(n6470), .C(wclk), .QN(n5100) );
  DFE1 \mem_reg_43][11  ( .D(D_11), .E(n6470), .C(wclk), .QN(n5101) );
  DFE1 \mem_reg_43][10  ( .D(D_10), .E(n6470), .C(wclk), .QN(n5102) );
  DFE1 \mem_reg_43][9  ( .D(D_9), .E(n6470), .C(wclk), .QN(n5103) );
  DFE1 \mem_reg_43][8  ( .D(D_8), .E(n6470), .C(wclk), .QN(n5104) );
  DFE1 \mem_reg_43][7  ( .D(D_7), .E(n6470), .C(wclk), .QN(n5105) );
  DFE1 \mem_reg_43][6  ( .D(D_6), .E(n6470), .C(wclk), .QN(n5106) );
  DFE1 \mem_reg_43][5  ( .D(D_5), .E(n6470), .C(wclk), .QN(n5107) );
  DFE1 \mem_reg_43][4  ( .D(D_4), .E(n6470), .C(wclk), .QN(n5108) );
  DFE1 \mem_reg_43][3  ( .D(D_3), .E(n6470), .C(wclk), .QN(n5109) );
  DFE1 \mem_reg_43][2  ( .D(D_2), .E(n6470), .C(wclk), .QN(n5110) );
  DFE1 \mem_reg_43][1  ( .D(D_1), .E(n6470), .C(wclk), .QN(n5111) );
  DFE1 \mem_reg_43][0  ( .D(D_0), .E(n6470), .C(wclk), .QN(n5112) );
  DFE1 \mem_reg_42][23  ( .D(D_23), .E(n6469), .C(wclk), .QN(n5113) );
  DFE1 \mem_reg_42][22  ( .D(D_22), .E(n6469), .C(wclk), .QN(n5114) );
  DFE1 \mem_reg_42][21  ( .D(D_21), .E(n6469), .C(wclk), .QN(n5115) );
  DFE1 \mem_reg_42][20  ( .D(D_20), .E(n6469), .C(wclk), .QN(n5116) );
  DFE1 \mem_reg_42][19  ( .D(D_19), .E(n6469), .C(wclk), .QN(n5117) );
  DFE1 \mem_reg_42][18  ( .D(D_18), .E(n6469), .C(wclk), .QN(n5118) );
  DFE1 \mem_reg_42][17  ( .D(D_17), .E(n6469), .C(wclk), .QN(n5119) );
  DFE1 \mem_reg_42][16  ( .D(D_16), .E(n6469), .C(wclk), .QN(n5120) );
  DFE1 \mem_reg_42][15  ( .D(D_15), .E(n6469), .C(wclk), .QN(n5121) );
  DFE1 \mem_reg_42][14  ( .D(D_14), .E(n6469), .C(wclk), .QN(n5122) );
  DFE1 \mem_reg_42][13  ( .D(D_13), .E(n6469), .C(wclk), .QN(n5123) );
  DFE1 \mem_reg_42][12  ( .D(D_12), .E(n6469), .C(wclk), .QN(n5124) );
  DFE1 \mem_reg_42][11  ( .D(D_11), .E(n6469), .C(wclk), .QN(n5125) );
  DFE1 \mem_reg_42][10  ( .D(D_10), .E(n6469), .C(wclk), .QN(n5126) );
  DFE1 \mem_reg_42][9  ( .D(D_9), .E(n6469), .C(wclk), .QN(n5127) );
  DFE1 \mem_reg_42][8  ( .D(D_8), .E(n6469), .C(wclk), .QN(n5128) );
  DFE1 \mem_reg_42][7  ( .D(D_7), .E(n6469), .C(wclk), .QN(n5129) );
  DFE1 \mem_reg_42][6  ( .D(D_6), .E(n6469), .C(wclk), .QN(n5130) );
  DFE1 \mem_reg_42][5  ( .D(D_5), .E(n6469), .C(wclk), .QN(n5131) );
  DFE1 \mem_reg_42][4  ( .D(D_4), .E(n6469), .C(wclk), .QN(n5132) );
  DFE1 \mem_reg_42][3  ( .D(D_3), .E(n6469), .C(wclk), .QN(n5133) );
  DFE1 \mem_reg_42][2  ( .D(D_2), .E(n6469), .C(wclk), .QN(n5134) );
  DFE1 \mem_reg_42][1  ( .D(D_1), .E(n6469), .C(wclk), .QN(n5135) );
  DFE1 \mem_reg_42][0  ( .D(D_0), .E(n6469), .C(wclk), .QN(n5136) );
  DFE1 \mem_reg_41][23  ( .D(D_23), .E(n6468), .C(wclk), .QN(n5137) );
  DFE1 \mem_reg_41][22  ( .D(D_22), .E(n6468), .C(wclk), .QN(n5138) );
  DFE1 \mem_reg_41][21  ( .D(D_21), .E(n6468), .C(wclk), .QN(n5139) );
  DFE1 \mem_reg_41][20  ( .D(D_20), .E(n6468), .C(wclk), .QN(n5140) );
  DFE1 \mem_reg_41][19  ( .D(D_19), .E(n6468), .C(wclk), .QN(n5141) );
  DFE1 \mem_reg_41][18  ( .D(D_18), .E(n6468), .C(wclk), .QN(n5142) );
  DFE1 \mem_reg_41][17  ( .D(D_17), .E(n6468), .C(wclk), .QN(n5143) );
  DFE1 \mem_reg_41][16  ( .D(D_16), .E(n6468), .C(wclk), .QN(n5144) );
  DFE1 \mem_reg_41][15  ( .D(D_15), .E(n6468), .C(wclk), .QN(n5145) );
  DFE1 \mem_reg_41][14  ( .D(D_14), .E(n6468), .C(wclk), .QN(n5146) );
  DFE1 \mem_reg_41][13  ( .D(D_13), .E(n6468), .C(wclk), .QN(n5147) );
  DFE1 \mem_reg_41][12  ( .D(D_12), .E(n6468), .C(wclk), .QN(n5148) );
  DFE1 \mem_reg_41][11  ( .D(D_11), .E(n6468), .C(wclk), .QN(n5149) );
  DFE1 \mem_reg_41][10  ( .D(D_10), .E(n6468), .C(wclk), .QN(n5150) );
  DFE1 \mem_reg_41][9  ( .D(D_9), .E(n6468), .C(wclk), .QN(n5151) );
  DFE1 \mem_reg_41][8  ( .D(D_8), .E(n6468), .C(wclk), .QN(n5152) );
  DFE1 \mem_reg_41][7  ( .D(D_7), .E(n6468), .C(wclk), .QN(n5153) );
  DFE1 \mem_reg_41][6  ( .D(D_6), .E(n6468), .C(wclk), .QN(n5154) );
  DFE1 \mem_reg_41][5  ( .D(D_5), .E(n6468), .C(wclk), .QN(n5155) );
  DFE1 \mem_reg_41][4  ( .D(D_4), .E(n6468), .C(wclk), .QN(n5156) );
  DFE1 \mem_reg_41][3  ( .D(D_3), .E(n6468), .C(wclk), .QN(n5157) );
  DFE1 \mem_reg_41][2  ( .D(D_2), .E(n6468), .C(wclk), .QN(n5158) );
  DFE1 \mem_reg_41][1  ( .D(D_1), .E(n6468), .C(wclk), .QN(n5159) );
  DFE1 \mem_reg_41][0  ( .D(D_0), .E(n6468), .C(wclk), .QN(n5160) );
  DFE1 \mem_reg_40][23  ( .D(D_23), .E(n6467), .C(wclk), .QN(n5161) );
  DFE1 \mem_reg_40][22  ( .D(D_22), .E(n6467), .C(wclk), .QN(n5162) );
  DFE1 \mem_reg_40][21  ( .D(D_21), .E(n6467), .C(wclk), .QN(n5163) );
  DFE1 \mem_reg_40][20  ( .D(D_20), .E(n6467), .C(wclk), .QN(n5164) );
  DFE1 \mem_reg_40][19  ( .D(D_19), .E(n6467), .C(wclk), .QN(n5165) );
  DFE1 \mem_reg_40][18  ( .D(D_18), .E(n6467), .C(wclk), .QN(n5166) );
  DFE1 \mem_reg_40][17  ( .D(D_17), .E(n6467), .C(wclk), .QN(n5167) );
  DFE1 \mem_reg_40][16  ( .D(D_16), .E(n6467), .C(wclk), .QN(n5168) );
  DFE1 \mem_reg_40][15  ( .D(D_15), .E(n6467), .C(wclk), .QN(n5169) );
  DFE1 \mem_reg_40][14  ( .D(D_14), .E(n6467), .C(wclk), .QN(n5170) );
  DFE1 \mem_reg_40][13  ( .D(D_13), .E(n6467), .C(wclk), .QN(n5171) );
  DFE1 \mem_reg_40][12  ( .D(D_12), .E(n6467), .C(wclk), .QN(n5172) );
  DFE1 \mem_reg_40][11  ( .D(D_11), .E(n6467), .C(wclk), .QN(n5173) );
  DFE1 \mem_reg_40][10  ( .D(D_10), .E(n6467), .C(wclk), .QN(n5174) );
  DFE1 \mem_reg_40][9  ( .D(D_9), .E(n6467), .C(wclk), .QN(n5175) );
  DFE1 \mem_reg_40][8  ( .D(D_8), .E(n6467), .C(wclk), .QN(n5176) );
  DFE1 \mem_reg_40][7  ( .D(D_7), .E(n6467), .C(wclk), .QN(n5177) );
  DFE1 \mem_reg_40][6  ( .D(D_6), .E(n6467), .C(wclk), .QN(n5178) );
  DFE1 \mem_reg_40][5  ( .D(D_5), .E(n6467), .C(wclk), .QN(n5179) );
  DFE1 \mem_reg_40][4  ( .D(D_4), .E(n6467), .C(wclk), .QN(n5180) );
  DFE1 \mem_reg_40][3  ( .D(D_3), .E(n6467), .C(wclk), .QN(n5181) );
  DFE1 \mem_reg_40][2  ( .D(D_2), .E(n6467), .C(wclk), .QN(n5182) );
  DFE1 \mem_reg_40][1  ( .D(D_1), .E(n6467), .C(wclk), .QN(n5183) );
  DFE1 \mem_reg_40][0  ( .D(D_0), .E(n6467), .C(wclk), .QN(n5184) );
  DFE1 \mem_reg_39][23  ( .D(D_23), .E(n6466), .C(wclk), .QN(n5185) );
  DFE1 \mem_reg_39][22  ( .D(D_22), .E(n6466), .C(wclk), .QN(n5186) );
  DFE1 \mem_reg_39][21  ( .D(D_21), .E(n6466), .C(wclk), .QN(n5187) );
  DFE1 \mem_reg_39][20  ( .D(D_20), .E(n6466), .C(wclk), .QN(n5188) );
  DFE1 \mem_reg_39][19  ( .D(D_19), .E(n6466), .C(wclk), .QN(n5189) );
  DFE1 \mem_reg_39][18  ( .D(D_18), .E(n6466), .C(wclk), .QN(n5190) );
  DFE1 \mem_reg_39][17  ( .D(D_17), .E(n6466), .C(wclk), .QN(n5191) );
  DFE1 \mem_reg_39][16  ( .D(D_16), .E(n6466), .C(wclk), .QN(n5192) );
  DFE1 \mem_reg_39][15  ( .D(D_15), .E(n6466), .C(wclk), .QN(n5193) );
  DFE1 \mem_reg_39][14  ( .D(D_14), .E(n6466), .C(wclk), .QN(n5194) );
  DFE1 \mem_reg_39][13  ( .D(D_13), .E(n6466), .C(wclk), .QN(n5195) );
  DFE1 \mem_reg_39][12  ( .D(D_12), .E(n6466), .C(wclk), .QN(n5196) );
  DFE1 \mem_reg_39][11  ( .D(D_11), .E(n6466), .C(wclk), .QN(n5197) );
  DFE1 \mem_reg_39][10  ( .D(D_10), .E(n6466), .C(wclk), .QN(n5198) );
  DFE1 \mem_reg_39][9  ( .D(D_9), .E(n6466), .C(wclk), .QN(n5199) );
  DFE1 \mem_reg_39][8  ( .D(D_8), .E(n6466), .C(wclk), .QN(n5200) );
  DFE1 \mem_reg_39][7  ( .D(D_7), .E(n6466), .C(wclk), .QN(n5201) );
  DFE1 \mem_reg_39][6  ( .D(D_6), .E(n6466), .C(wclk), .QN(n5202) );
  DFE1 \mem_reg_39][5  ( .D(D_5), .E(n6466), .C(wclk), .QN(n5203) );
  DFE1 \mem_reg_39][4  ( .D(D_4), .E(n6466), .C(wclk), .QN(n5204) );
  DFE1 \mem_reg_39][3  ( .D(D_3), .E(n6466), .C(wclk), .QN(n5205) );
  DFE1 \mem_reg_39][2  ( .D(D_2), .E(n6466), .C(wclk), .QN(n5206) );
  DFE1 \mem_reg_39][1  ( .D(D_1), .E(n6466), .C(wclk), .QN(n5207) );
  DFE1 \mem_reg_39][0  ( .D(D_0), .E(n6466), .C(wclk), .QN(n5208) );
  DFE1 \mem_reg_38][23  ( .D(D_23), .E(n6465), .C(wclk), .QN(n5209) );
  DFE1 \mem_reg_38][22  ( .D(D_22), .E(n6465), .C(wclk), .QN(n5210) );
  DFE1 \mem_reg_38][21  ( .D(D_21), .E(n6465), .C(wclk), .QN(n5211) );
  DFE1 \mem_reg_38][20  ( .D(D_20), .E(n6465), .C(wclk), .QN(n5212) );
  DFE1 \mem_reg_38][19  ( .D(D_19), .E(n6465), .C(wclk), .QN(n5213) );
  DFE1 \mem_reg_38][18  ( .D(D_18), .E(n6465), .C(wclk), .QN(n5214) );
  DFE1 \mem_reg_38][17  ( .D(D_17), .E(n6465), .C(wclk), .QN(n5215) );
  DFE1 \mem_reg_38][16  ( .D(D_16), .E(n6465), .C(wclk), .QN(n5216) );
  DFE1 \mem_reg_38][15  ( .D(D_15), .E(n6465), .C(wclk), .QN(n5217) );
  DFE1 \mem_reg_38][14  ( .D(D_14), .E(n6465), .C(wclk), .QN(n5218) );
  DFE1 \mem_reg_38][13  ( .D(D_13), .E(n6465), .C(wclk), .QN(n5219) );
  DFE1 \mem_reg_38][12  ( .D(D_12), .E(n6465), .C(wclk), .QN(n5220) );
  DFE1 \mem_reg_38][11  ( .D(D_11), .E(n6465), .C(wclk), .QN(n5221) );
  DFE1 \mem_reg_38][10  ( .D(D_10), .E(n6465), .C(wclk), .QN(n5222) );
  DFE1 \mem_reg_38][9  ( .D(D_9), .E(n6465), .C(wclk), .QN(n5223) );
  DFE1 \mem_reg_38][8  ( .D(D_8), .E(n6465), .C(wclk), .QN(n5224) );
  DFE1 \mem_reg_38][7  ( .D(D_7), .E(n6465), .C(wclk), .QN(n5225) );
  DFE1 \mem_reg_38][6  ( .D(D_6), .E(n6465), .C(wclk), .QN(n5226) );
  DFE1 \mem_reg_38][5  ( .D(D_5), .E(n6465), .C(wclk), .QN(n5227) );
  DFE1 \mem_reg_38][4  ( .D(D_4), .E(n6465), .C(wclk), .QN(n5228) );
  DFE1 \mem_reg_38][3  ( .D(D_3), .E(n6465), .C(wclk), .QN(n5229) );
  DFE1 \mem_reg_38][2  ( .D(D_2), .E(n6465), .C(wclk), .QN(n5230) );
  DFE1 \mem_reg_38][1  ( .D(D_1), .E(n6465), .C(wclk), .QN(n5231) );
  DFE1 \mem_reg_38][0  ( .D(D_0), .E(n6465), .C(wclk), .QN(n5232) );
  DFE1 \mem_reg_37][23  ( .D(D_23), .E(n6464), .C(wclk), .QN(n5233) );
  DFE1 \mem_reg_37][22  ( .D(D_22), .E(n6464), .C(wclk), .QN(n5234) );
  DFE1 \mem_reg_37][21  ( .D(D_21), .E(n6464), .C(wclk), .QN(n5235) );
  DFE1 \mem_reg_37][20  ( .D(D_20), .E(n6464), .C(wclk), .QN(n5236) );
  DFE1 \mem_reg_37][19  ( .D(D_19), .E(n6464), .C(wclk), .QN(n5237) );
  DFE1 \mem_reg_37][18  ( .D(D_18), .E(n6464), .C(wclk), .QN(n5238) );
  DFE1 \mem_reg_37][17  ( .D(D_17), .E(n6464), .C(wclk), .QN(n5239) );
  DFE1 \mem_reg_37][16  ( .D(D_16), .E(n6464), .C(wclk), .QN(n5240) );
  DFE1 \mem_reg_37][15  ( .D(D_15), .E(n6464), .C(wclk), .QN(n5241) );
  DFE1 \mem_reg_37][14  ( .D(D_14), .E(n6464), .C(wclk), .QN(n5242) );
  DFE1 \mem_reg_37][13  ( .D(D_13), .E(n6464), .C(wclk), .QN(n5243) );
  DFE1 \mem_reg_37][12  ( .D(D_12), .E(n6464), .C(wclk), .QN(n5244) );
  DFE1 \mem_reg_37][11  ( .D(D_11), .E(n6464), .C(wclk), .QN(n5245) );
  DFE1 \mem_reg_37][10  ( .D(D_10), .E(n6464), .C(wclk), .QN(n5246) );
  DFE1 \mem_reg_37][9  ( .D(D_9), .E(n6464), .C(wclk), .QN(n5247) );
  DFE1 \mem_reg_37][8  ( .D(D_8), .E(n6464), .C(wclk), .QN(n5248) );
  DFE1 \mem_reg_37][7  ( .D(D_7), .E(n6464), .C(wclk), .QN(n5249) );
  DFE1 \mem_reg_37][6  ( .D(D_6), .E(n6464), .C(wclk), .QN(n5250) );
  DFE1 \mem_reg_37][5  ( .D(D_5), .E(n6464), .C(wclk), .QN(n5251) );
  DFE1 \mem_reg_37][4  ( .D(D_4), .E(n6464), .C(wclk), .QN(n5252) );
  DFE1 \mem_reg_37][3  ( .D(D_3), .E(n6464), .C(wclk), .QN(n5253) );
  DFE1 \mem_reg_37][2  ( .D(D_2), .E(n6464), .C(wclk), .QN(n5254) );
  DFE1 \mem_reg_37][1  ( .D(D_1), .E(n6464), .C(wclk), .QN(n5255) );
  DFE1 \mem_reg_37][0  ( .D(D_0), .E(n6464), .C(wclk), .QN(n5256) );
  DFE1 \mem_reg_36][23  ( .D(D_23), .E(n6463), .C(wclk), .QN(n5257) );
  DFE1 \mem_reg_36][22  ( .D(D_22), .E(n6463), .C(wclk), .QN(n5258) );
  DFE1 \mem_reg_36][21  ( .D(D_21), .E(n6463), .C(wclk), .QN(n5259) );
  DFE1 \mem_reg_36][20  ( .D(D_20), .E(n6463), .C(wclk), .QN(n5260) );
  DFE1 \mem_reg_36][19  ( .D(D_19), .E(n6463), .C(wclk), .QN(n5261) );
  DFE1 \mem_reg_36][18  ( .D(D_18), .E(n6463), .C(wclk), .QN(n5262) );
  DFE1 \mem_reg_36][17  ( .D(D_17), .E(n6463), .C(wclk), .QN(n5263) );
  DFE1 \mem_reg_36][16  ( .D(D_16), .E(n6463), .C(wclk), .QN(n5264) );
  DFE1 \mem_reg_36][15  ( .D(D_15), .E(n6463), .C(wclk), .QN(n5265) );
  DFE1 \mem_reg_36][14  ( .D(D_14), .E(n6463), .C(wclk), .QN(n5266) );
  DFE1 \mem_reg_36][13  ( .D(D_13), .E(n6463), .C(wclk), .QN(n5267) );
  DFE1 \mem_reg_36][12  ( .D(D_12), .E(n6463), .C(wclk), .QN(n5268) );
  DFE1 \mem_reg_36][11  ( .D(D_11), .E(n6463), .C(wclk), .QN(n5269) );
  DFE1 \mem_reg_36][10  ( .D(D_10), .E(n6463), .C(wclk), .QN(n5270) );
  DFE1 \mem_reg_36][9  ( .D(D_9), .E(n6463), .C(wclk), .QN(n5271) );
  DFE1 \mem_reg_36][8  ( .D(D_8), .E(n6463), .C(wclk), .QN(n5272) );
  DFE1 \mem_reg_36][7  ( .D(D_7), .E(n6463), .C(wclk), .QN(n5273) );
  DFE1 \mem_reg_36][6  ( .D(D_6), .E(n6463), .C(wclk), .QN(n5274) );
  DFE1 \mem_reg_36][5  ( .D(D_5), .E(n6463), .C(wclk), .QN(n5275) );
  DFE1 \mem_reg_36][4  ( .D(D_4), .E(n6463), .C(wclk), .QN(n5276) );
  DFE1 \mem_reg_36][3  ( .D(D_3), .E(n6463), .C(wclk), .QN(n5277) );
  DFE1 \mem_reg_36][2  ( .D(D_2), .E(n6463), .C(wclk), .QN(n5278) );
  DFE1 \mem_reg_36][1  ( .D(D_1), .E(n6463), .C(wclk), .QN(n5279) );
  DFE1 \mem_reg_36][0  ( .D(D_0), .E(n6463), .C(wclk), .QN(n5280) );
  DFE1 \mem_reg_35][23  ( .D(D_23), .E(n6462), .C(wclk), .QN(n5281) );
  DFE1 \mem_reg_35][22  ( .D(D_22), .E(n6462), .C(wclk), .QN(n5282) );
  DFE1 \mem_reg_35][21  ( .D(D_21), .E(n6462), .C(wclk), .QN(n5283) );
  DFE1 \mem_reg_35][20  ( .D(D_20), .E(n6462), .C(wclk), .QN(n5284) );
  DFE1 \mem_reg_35][19  ( .D(D_19), .E(n6462), .C(wclk), .QN(n5285) );
  DFE1 \mem_reg_35][18  ( .D(D_18), .E(n6462), .C(wclk), .QN(n5286) );
  DFE1 \mem_reg_35][17  ( .D(D_17), .E(n6462), .C(wclk), .QN(n5287) );
  DFE1 \mem_reg_35][16  ( .D(D_16), .E(n6462), .C(wclk), .QN(n5288) );
  DFE1 \mem_reg_35][15  ( .D(D_15), .E(n6462), .C(wclk), .QN(n5289) );
  DFE1 \mem_reg_35][14  ( .D(D_14), .E(n6462), .C(wclk), .QN(n5290) );
  DFE1 \mem_reg_35][13  ( .D(D_13), .E(n6462), .C(wclk), .QN(n5291) );
  DFE1 \mem_reg_35][12  ( .D(D_12), .E(n6462), .C(wclk), .QN(n5292) );
  DFE1 \mem_reg_35][11  ( .D(D_11), .E(n6462), .C(wclk), .QN(n5293) );
  DFE1 \mem_reg_35][10  ( .D(D_10), .E(n6462), .C(wclk), .QN(n5294) );
  DFE1 \mem_reg_35][9  ( .D(D_9), .E(n6462), .C(wclk), .QN(n5295) );
  DFE1 \mem_reg_35][8  ( .D(D_8), .E(n6462), .C(wclk), .QN(n5296) );
  DFE1 \mem_reg_35][7  ( .D(D_7), .E(n6462), .C(wclk), .QN(n5297) );
  DFE1 \mem_reg_35][6  ( .D(D_6), .E(n6462), .C(wclk), .QN(n5298) );
  DFE1 \mem_reg_35][5  ( .D(D_5), .E(n6462), .C(wclk), .QN(n5299) );
  DFE1 \mem_reg_35][4  ( .D(D_4), .E(n6462), .C(wclk), .QN(n5300) );
  DFE1 \mem_reg_35][3  ( .D(D_3), .E(n6462), .C(wclk), .QN(n5301) );
  DFE1 \mem_reg_35][2  ( .D(D_2), .E(n6462), .C(wclk), .QN(n5302) );
  DFE1 \mem_reg_35][1  ( .D(D_1), .E(n6462), .C(wclk), .QN(n5303) );
  DFE1 \mem_reg_35][0  ( .D(D_0), .E(n6462), .C(wclk), .QN(n5304) );
  DFE1 \mem_reg_34][23  ( .D(D_23), .E(n6461), .C(wclk), .QN(n5305) );
  DFE1 \mem_reg_34][22  ( .D(D_22), .E(n6461), .C(wclk), .QN(n5306) );
  DFE1 \mem_reg_34][21  ( .D(D_21), .E(n6461), .C(wclk), .QN(n5307) );
  DFE1 \mem_reg_34][20  ( .D(D_20), .E(n6461), .C(wclk), .QN(n5308) );
  DFE1 \mem_reg_34][19  ( .D(D_19), .E(n6461), .C(wclk), .QN(n5309) );
  DFE1 \mem_reg_34][18  ( .D(D_18), .E(n6461), .C(wclk), .QN(n5310) );
  DFE1 \mem_reg_34][17  ( .D(D_17), .E(n6461), .C(wclk), .QN(n5311) );
  DFE1 \mem_reg_34][16  ( .D(D_16), .E(n6461), .C(wclk), .QN(n5312) );
  DFE1 \mem_reg_34][15  ( .D(D_15), .E(n6461), .C(wclk), .QN(n5313) );
  DFE1 \mem_reg_34][14  ( .D(D_14), .E(n6461), .C(wclk), .QN(n5314) );
  DFE1 \mem_reg_34][13  ( .D(D_13), .E(n6461), .C(wclk), .QN(n5315) );
  DFE1 \mem_reg_34][12  ( .D(D_12), .E(n6461), .C(wclk), .QN(n5316) );
  DFE1 \mem_reg_34][11  ( .D(D_11), .E(n6461), .C(wclk), .QN(n5317) );
  DFE1 \mem_reg_34][10  ( .D(D_10), .E(n6461), .C(wclk), .QN(n5318) );
  DFE1 \mem_reg_34][9  ( .D(D_9), .E(n6461), .C(wclk), .QN(n5319) );
  DFE1 \mem_reg_34][8  ( .D(D_8), .E(n6461), .C(wclk), .QN(n5320) );
  DFE1 \mem_reg_34][7  ( .D(D_7), .E(n6461), .C(wclk), .QN(n5321) );
  DFE1 \mem_reg_34][6  ( .D(D_6), .E(n6461), .C(wclk), .QN(n5322) );
  DFE1 \mem_reg_34][5  ( .D(D_5), .E(n6461), .C(wclk), .QN(n5323) );
  DFE1 \mem_reg_34][4  ( .D(D_4), .E(n6461), .C(wclk), .QN(n5324) );
  DFE1 \mem_reg_34][3  ( .D(D_3), .E(n6461), .C(wclk), .QN(n5325) );
  DFE1 \mem_reg_34][2  ( .D(D_2), .E(n6461), .C(wclk), .QN(n5326) );
  DFE1 \mem_reg_34][1  ( .D(D_1), .E(n6461), .C(wclk), .QN(n5327) );
  DFE1 \mem_reg_34][0  ( .D(D_0), .E(n6461), .C(wclk), .QN(n5328) );
  DFE1 \mem_reg_33][23  ( .D(D_23), .E(n6459), .C(wclk), .QN(n5329) );
  DFE1 \mem_reg_33][22  ( .D(D_22), .E(n6459), .C(wclk), .QN(n5330) );
  DFE1 \mem_reg_33][21  ( .D(D_21), .E(n6459), .C(wclk), .QN(n5331) );
  DFE1 \mem_reg_33][20  ( .D(D_20), .E(n6459), .C(wclk), .QN(n5332) );
  DFE1 \mem_reg_33][19  ( .D(D_19), .E(n6459), .C(wclk), .QN(n5333) );
  DFE1 \mem_reg_33][18  ( .D(D_18), .E(n6459), .C(wclk), .QN(n5334) );
  DFE1 \mem_reg_33][17  ( .D(D_17), .E(n6459), .C(wclk), .QN(n5335) );
  DFE1 \mem_reg_33][16  ( .D(D_16), .E(n6459), .C(wclk), .QN(n5336) );
  DFE1 \mem_reg_33][15  ( .D(D_15), .E(n6459), .C(wclk), .QN(n5337) );
  DFE1 \mem_reg_33][14  ( .D(D_14), .E(n6459), .C(wclk), .QN(n5338) );
  DFE1 \mem_reg_33][13  ( .D(D_13), .E(n6459), .C(wclk), .QN(n5339) );
  DFE1 \mem_reg_33][12  ( .D(D_12), .E(n6459), .C(wclk), .QN(n5340) );
  DFE1 \mem_reg_33][11  ( .D(D_11), .E(n6459), .C(wclk), .QN(n5341) );
  DFE1 \mem_reg_33][10  ( .D(D_10), .E(n6459), .C(wclk), .QN(n5342) );
  DFE1 \mem_reg_33][9  ( .D(D_9), .E(n6459), .C(wclk), .QN(n5343) );
  DFE1 \mem_reg_33][8  ( .D(D_8), .E(n6459), .C(wclk), .QN(n5344) );
  DFE1 \mem_reg_33][7  ( .D(D_7), .E(n6459), .C(wclk), .QN(n5345) );
  DFE1 \mem_reg_33][6  ( .D(D_6), .E(n6459), .C(wclk), .QN(n5346) );
  DFE1 \mem_reg_33][5  ( .D(D_5), .E(n6459), .C(wclk), .QN(n5347) );
  DFE1 \mem_reg_33][4  ( .D(D_4), .E(n6459), .C(wclk), .QN(n5348) );
  DFE1 \mem_reg_33][3  ( .D(D_3), .E(n6459), .C(wclk), .QN(n5349) );
  DFE1 \mem_reg_33][2  ( .D(D_2), .E(n6459), .C(wclk), .QN(n5350) );
  DFE1 \mem_reg_33][1  ( .D(D_1), .E(n6459), .C(wclk), .QN(n5351) );
  DFE1 \mem_reg_33][0  ( .D(D_0), .E(n6459), .C(wclk), .QN(n5352) );
  DFE1 \mem_reg_32][23  ( .D(D_23), .E(n6457), .C(wclk), .QN(n5353) );
  DFE1 \mem_reg_32][22  ( .D(D_22), .E(n6457), .C(wclk), .QN(n5354) );
  DFE1 \mem_reg_32][21  ( .D(D_21), .E(n6457), .C(wclk), .QN(n5355) );
  DFE1 \mem_reg_32][20  ( .D(D_20), .E(n6457), .C(wclk), .QN(n5356) );
  DFE1 \mem_reg_32][19  ( .D(D_19), .E(n6457), .C(wclk), .QN(n5357) );
  DFE1 \mem_reg_32][18  ( .D(D_18), .E(n6457), .C(wclk), .QN(n5358) );
  DFE1 \mem_reg_32][17  ( .D(D_17), .E(n6457), .C(wclk), .QN(n5359) );
  DFE1 \mem_reg_32][16  ( .D(D_16), .E(n6457), .C(wclk), .QN(n5360) );
  DFE1 \mem_reg_32][15  ( .D(D_15), .E(n6457), .C(wclk), .QN(n5361) );
  DFE1 \mem_reg_32][14  ( .D(D_14), .E(n6457), .C(wclk), .QN(n5362) );
  DFE1 \mem_reg_32][13  ( .D(D_13), .E(n6457), .C(wclk), .QN(n5363) );
  DFE1 \mem_reg_32][12  ( .D(D_12), .E(n6457), .C(wclk), .QN(n5364) );
  DFE1 \mem_reg_32][11  ( .D(D_11), .E(n6457), .C(wclk), .QN(n5365) );
  DFE1 \mem_reg_32][10  ( .D(D_10), .E(n6457), .C(wclk), .QN(n5366) );
  DFE1 \mem_reg_32][9  ( .D(D_9), .E(n6457), .C(wclk), .QN(n5367) );
  DFE1 \mem_reg_32][8  ( .D(D_8), .E(n6457), .C(wclk), .QN(n5368) );
  DFE1 \mem_reg_32][7  ( .D(D_7), .E(n6457), .C(wclk), .QN(n5369) );
  DFE1 \mem_reg_32][6  ( .D(D_6), .E(n6457), .C(wclk), .QN(n5370) );
  DFE1 \mem_reg_32][5  ( .D(D_5), .E(n6457), .C(wclk), .QN(n5371) );
  DFE1 \mem_reg_32][4  ( .D(D_4), .E(n6457), .C(wclk), .QN(n5372) );
  DFE1 \mem_reg_32][3  ( .D(D_3), .E(n6457), .C(wclk), .QN(n5373) );
  DFE1 \mem_reg_32][2  ( .D(D_2), .E(n6457), .C(wclk), .QN(n5374) );
  DFE1 \mem_reg_32][1  ( .D(D_1), .E(n6457), .C(wclk), .QN(n5375) );
  DFE1 \mem_reg_32][0  ( .D(D_0), .E(n6457), .C(wclk), .QN(n5376) );
  DFE1 \mem_reg_31][23  ( .D(D_23), .E(n6456), .C(wclk), .QN(n5377) );
  DFE1 \mem_reg_31][22  ( .D(D_22), .E(n6456), .C(wclk), .QN(n5378) );
  DFE1 \mem_reg_31][21  ( .D(D_21), .E(n6456), .C(wclk), .QN(n5379) );
  DFE1 \mem_reg_31][20  ( .D(D_20), .E(n6456), .C(wclk), .QN(n5380) );
  DFE1 \mem_reg_31][19  ( .D(D_19), .E(n6456), .C(wclk), .QN(n5381) );
  DFE1 \mem_reg_31][18  ( .D(D_18), .E(n6456), .C(wclk), .QN(n5382) );
  DFE1 \mem_reg_31][17  ( .D(D_17), .E(n6456), .C(wclk), .QN(n5383) );
  DFE1 \mem_reg_31][16  ( .D(D_16), .E(n6456), .C(wclk), .QN(n5384) );
  DFE1 \mem_reg_31][15  ( .D(D_15), .E(n6456), .C(wclk), .QN(n5385) );
  DFE1 \mem_reg_31][14  ( .D(D_14), .E(n6456), .C(wclk), .QN(n5386) );
  DFE1 \mem_reg_31][13  ( .D(D_13), .E(n6456), .C(wclk), .QN(n5387) );
  DFE1 \mem_reg_31][12  ( .D(D_12), .E(n6456), .C(wclk), .QN(n5388) );
  DFE1 \mem_reg_31][11  ( .D(D_11), .E(n6456), .C(wclk), .QN(n5389) );
  DFE1 \mem_reg_31][10  ( .D(D_10), .E(n6456), .C(wclk), .QN(n5390) );
  DFE1 \mem_reg_31][9  ( .D(D_9), .E(n6456), .C(wclk), .QN(n5391) );
  DFE1 \mem_reg_31][8  ( .D(D_8), .E(n6456), .C(wclk), .QN(n5392) );
  DFE1 \mem_reg_31][7  ( .D(D_7), .E(n6456), .C(wclk), .QN(n5393) );
  DFE1 \mem_reg_31][6  ( .D(D_6), .E(n6456), .C(wclk), .QN(n5394) );
  DFE1 \mem_reg_31][5  ( .D(D_5), .E(n6456), .C(wclk), .QN(n5395) );
  DFE1 \mem_reg_31][4  ( .D(D_4), .E(n6456), .C(wclk), .QN(n5396) );
  DFE1 \mem_reg_31][3  ( .D(D_3), .E(n6456), .C(wclk), .QN(n5397) );
  DFE1 \mem_reg_31][2  ( .D(D_2), .E(n6456), .C(wclk), .QN(n5398) );
  DFE1 \mem_reg_31][1  ( .D(D_1), .E(n6456), .C(wclk), .QN(n5399) );
  DFE1 \mem_reg_31][0  ( .D(D_0), .E(n6456), .C(wclk), .QN(n5400) );
  DFE1 \mem_reg_30][23  ( .D(D_23), .E(n6455), .C(wclk), .QN(n5401) );
  DFE1 \mem_reg_30][22  ( .D(D_22), .E(n6455), .C(wclk), .QN(n5402) );
  DFE1 \mem_reg_30][21  ( .D(D_21), .E(n6455), .C(wclk), .QN(n5403) );
  DFE1 \mem_reg_30][20  ( .D(D_20), .E(n6455), .C(wclk), .QN(n5404) );
  DFE1 \mem_reg_30][19  ( .D(D_19), .E(n6455), .C(wclk), .QN(n5405) );
  DFE1 \mem_reg_30][18  ( .D(D_18), .E(n6455), .C(wclk), .QN(n5406) );
  DFE1 \mem_reg_30][17  ( .D(D_17), .E(n6455), .C(wclk), .QN(n5407) );
  DFE1 \mem_reg_30][16  ( .D(D_16), .E(n6455), .C(wclk), .QN(n5408) );
  DFE1 \mem_reg_30][15  ( .D(D_15), .E(n6455), .C(wclk), .QN(n5409) );
  DFE1 \mem_reg_30][14  ( .D(D_14), .E(n6455), .C(wclk), .QN(n5410) );
  DFE1 \mem_reg_30][13  ( .D(D_13), .E(n6455), .C(wclk), .QN(n5411) );
  DFE1 \mem_reg_30][12  ( .D(D_12), .E(n6455), .C(wclk), .QN(n5412) );
  DFE1 \mem_reg_30][11  ( .D(D_11), .E(n6455), .C(wclk), .QN(n5413) );
  DFE1 \mem_reg_30][10  ( .D(D_10), .E(n6455), .C(wclk), .QN(n5414) );
  DFE1 \mem_reg_30][9  ( .D(D_9), .E(n6455), .C(wclk), .QN(n5415) );
  DFE1 \mem_reg_30][8  ( .D(D_8), .E(n6455), .C(wclk), .QN(n5416) );
  DFE1 \mem_reg_30][7  ( .D(D_7), .E(n6455), .C(wclk), .QN(n5417) );
  DFE1 \mem_reg_30][6  ( .D(D_6), .E(n6455), .C(wclk), .QN(n5418) );
  DFE1 \mem_reg_30][5  ( .D(D_5), .E(n6455), .C(wclk), .QN(n5419) );
  DFE1 \mem_reg_30][4  ( .D(D_4), .E(n6455), .C(wclk), .QN(n5420) );
  DFE1 \mem_reg_30][3  ( .D(D_3), .E(n6455), .C(wclk), .QN(n5421) );
  DFE1 \mem_reg_30][2  ( .D(D_2), .E(n6455), .C(wclk), .QN(n5422) );
  DFE1 \mem_reg_30][1  ( .D(D_1), .E(n6455), .C(wclk), .QN(n5423) );
  DFE1 \mem_reg_30][0  ( .D(D_0), .E(n6455), .C(wclk), .QN(n5424) );
  DFE1 \mem_reg_29][23  ( .D(D_23), .E(n6454), .C(wclk), .QN(n5425) );
  DFE1 \mem_reg_29][22  ( .D(D_22), .E(n6454), .C(wclk), .QN(n5426) );
  DFE1 \mem_reg_29][21  ( .D(D_21), .E(n6454), .C(wclk), .QN(n5427) );
  DFE1 \mem_reg_29][20  ( .D(D_20), .E(n6454), .C(wclk), .QN(n5428) );
  DFE1 \mem_reg_29][19  ( .D(D_19), .E(n6454), .C(wclk), .QN(n5429) );
  DFE1 \mem_reg_29][18  ( .D(D_18), .E(n6454), .C(wclk), .QN(n5430) );
  DFE1 \mem_reg_29][17  ( .D(D_17), .E(n6454), .C(wclk), .QN(n5431) );
  DFE1 \mem_reg_29][16  ( .D(D_16), .E(n6454), .C(wclk), .QN(n5432) );
  DFE1 \mem_reg_29][15  ( .D(D_15), .E(n6454), .C(wclk), .QN(n5433) );
  DFE1 \mem_reg_29][14  ( .D(D_14), .E(n6454), .C(wclk), .QN(n5434) );
  DFE1 \mem_reg_29][13  ( .D(D_13), .E(n6454), .C(wclk), .QN(n5435) );
  DFE1 \mem_reg_29][12  ( .D(D_12), .E(n6454), .C(wclk), .QN(n5436) );
  DFE1 \mem_reg_29][11  ( .D(D_11), .E(n6454), .C(wclk), .QN(n5437) );
  DFE1 \mem_reg_29][10  ( .D(D_10), .E(n6454), .C(wclk), .QN(n5438) );
  DFE1 \mem_reg_29][9  ( .D(D_9), .E(n6454), .C(wclk), .QN(n5439) );
  DFE1 \mem_reg_29][8  ( .D(D_8), .E(n6454), .C(wclk), .QN(n5440) );
  DFE1 \mem_reg_29][7  ( .D(D_7), .E(n6454), .C(wclk), .QN(n5441) );
  DFE1 \mem_reg_29][6  ( .D(D_6), .E(n6454), .C(wclk), .QN(n5442) );
  DFE1 \mem_reg_29][5  ( .D(D_5), .E(n6454), .C(wclk), .QN(n5443) );
  DFE1 \mem_reg_29][4  ( .D(D_4), .E(n6454), .C(wclk), .QN(n5444) );
  DFE1 \mem_reg_29][3  ( .D(D_3), .E(n6454), .C(wclk), .QN(n5445) );
  DFE1 \mem_reg_29][2  ( .D(D_2), .E(n6454), .C(wclk), .QN(n5446) );
  DFE1 \mem_reg_29][1  ( .D(D_1), .E(n6454), .C(wclk), .QN(n5447) );
  DFE1 \mem_reg_29][0  ( .D(D_0), .E(n6454), .C(wclk), .QN(n5448) );
  DFE1 \mem_reg_28][23  ( .D(D_23), .E(n6453), .C(wclk), .QN(n5449) );
  DFE1 \mem_reg_28][22  ( .D(D_22), .E(n6453), .C(wclk), .QN(n5450) );
  DFE1 \mem_reg_28][21  ( .D(D_21), .E(n6453), .C(wclk), .QN(n5451) );
  DFE1 \mem_reg_28][20  ( .D(D_20), .E(n6453), .C(wclk), .QN(n5452) );
  DFE1 \mem_reg_28][19  ( .D(D_19), .E(n6453), .C(wclk), .QN(n5453) );
  DFE1 \mem_reg_28][18  ( .D(D_18), .E(n6453), .C(wclk), .QN(n5454) );
  DFE1 \mem_reg_28][17  ( .D(D_17), .E(n6453), .C(wclk), .QN(n5455) );
  DFE1 \mem_reg_28][16  ( .D(D_16), .E(n6453), .C(wclk), .QN(n5456) );
  DFE1 \mem_reg_28][15  ( .D(D_15), .E(n6453), .C(wclk), .QN(n5457) );
  DFE1 \mem_reg_28][14  ( .D(D_14), .E(n6453), .C(wclk), .QN(n5458) );
  DFE1 \mem_reg_28][13  ( .D(D_13), .E(n6453), .C(wclk), .QN(n5459) );
  DFE1 \mem_reg_28][12  ( .D(D_12), .E(n6453), .C(wclk), .QN(n5460) );
  DFE1 \mem_reg_28][11  ( .D(D_11), .E(n6453), .C(wclk), .QN(n5461) );
  DFE1 \mem_reg_28][10  ( .D(D_10), .E(n6453), .C(wclk), .QN(n5462) );
  DFE1 \mem_reg_28][9  ( .D(D_9), .E(n6453), .C(wclk), .QN(n5463) );
  DFE1 \mem_reg_28][8  ( .D(D_8), .E(n6453), .C(wclk), .QN(n5464) );
  DFE1 \mem_reg_28][7  ( .D(D_7), .E(n6453), .C(wclk), .QN(n5465) );
  DFE1 \mem_reg_28][6  ( .D(D_6), .E(n6453), .C(wclk), .QN(n5466) );
  DFE1 \mem_reg_28][5  ( .D(D_5), .E(n6453), .C(wclk), .QN(n5467) );
  DFE1 \mem_reg_28][4  ( .D(D_4), .E(n6453), .C(wclk), .QN(n5468) );
  DFE1 \mem_reg_28][3  ( .D(D_3), .E(n6453), .C(wclk), .QN(n5469) );
  DFE1 \mem_reg_28][2  ( .D(D_2), .E(n6453), .C(wclk), .QN(n5470) );
  DFE1 \mem_reg_28][1  ( .D(D_1), .E(n6453), .C(wclk), .QN(n5471) );
  DFE1 \mem_reg_28][0  ( .D(D_0), .E(n6453), .C(wclk), .QN(n5472) );
  DFE1 \mem_reg_27][23  ( .D(D_23), .E(n6452), .C(wclk), .QN(n5473) );
  DFE1 \mem_reg_27][22  ( .D(D_22), .E(n6452), .C(wclk), .QN(n5474) );
  DFE1 \mem_reg_27][21  ( .D(D_21), .E(n6452), .C(wclk), .QN(n5475) );
  DFE1 \mem_reg_27][20  ( .D(D_20), .E(n6452), .C(wclk), .QN(n5476) );
  DFE1 \mem_reg_27][19  ( .D(D_19), .E(n6452), .C(wclk), .QN(n5477) );
  DFE1 \mem_reg_27][18  ( .D(D_18), .E(n6452), .C(wclk), .QN(n5478) );
  DFE1 \mem_reg_27][17  ( .D(D_17), .E(n6452), .C(wclk), .QN(n5479) );
  DFE1 \mem_reg_27][16  ( .D(D_16), .E(n6452), .C(wclk), .QN(n5480) );
  DFE1 \mem_reg_27][15  ( .D(D_15), .E(n6452), .C(wclk), .QN(n5481) );
  DFE1 \mem_reg_27][14  ( .D(D_14), .E(n6452), .C(wclk), .QN(n5482) );
  DFE1 \mem_reg_27][13  ( .D(D_13), .E(n6452), .C(wclk), .QN(n5483) );
  DFE1 \mem_reg_27][12  ( .D(D_12), .E(n6452), .C(wclk), .QN(n5484) );
  DFE1 \mem_reg_27][11  ( .D(D_11), .E(n6452), .C(wclk), .QN(n5485) );
  DFE1 \mem_reg_27][10  ( .D(D_10), .E(n6452), .C(wclk), .QN(n5486) );
  DFE1 \mem_reg_27][9  ( .D(D_9), .E(n6452), .C(wclk), .QN(n5487) );
  DFE1 \mem_reg_27][8  ( .D(D_8), .E(n6452), .C(wclk), .QN(n5488) );
  DFE1 \mem_reg_27][7  ( .D(D_7), .E(n6452), .C(wclk), .QN(n5489) );
  DFE1 \mem_reg_27][6  ( .D(D_6), .E(n6452), .C(wclk), .QN(n5490) );
  DFE1 \mem_reg_27][5  ( .D(D_5), .E(n6452), .C(wclk), .QN(n5491) );
  DFE1 \mem_reg_27][4  ( .D(D_4), .E(n6452), .C(wclk), .QN(n5492) );
  DFE1 \mem_reg_27][3  ( .D(D_3), .E(n6452), .C(wclk), .QN(n5493) );
  DFE1 \mem_reg_27][2  ( .D(D_2), .E(n6452), .C(wclk), .QN(n5494) );
  DFE1 \mem_reg_27][1  ( .D(D_1), .E(n6452), .C(wclk), .QN(n5495) );
  DFE1 \mem_reg_27][0  ( .D(D_0), .E(n6452), .C(wclk), .QN(n5496) );
  DFE1 \mem_reg_26][23  ( .D(D_23), .E(n6451), .C(wclk), .QN(n5497) );
  DFE1 \mem_reg_26][22  ( .D(D_22), .E(n6451), .C(wclk), .QN(n5498) );
  DFE1 \mem_reg_26][21  ( .D(D_21), .E(n6451), .C(wclk), .QN(n5499) );
  DFE1 \mem_reg_26][20  ( .D(D_20), .E(n6451), .C(wclk), .QN(n5500) );
  DFE1 \mem_reg_26][19  ( .D(D_19), .E(n6451), .C(wclk), .QN(n5501) );
  DFE1 \mem_reg_26][18  ( .D(D_18), .E(n6451), .C(wclk), .QN(n5502) );
  DFE1 \mem_reg_26][17  ( .D(D_17), .E(n6451), .C(wclk), .QN(n5503) );
  DFE1 \mem_reg_26][16  ( .D(D_16), .E(n6451), .C(wclk), .QN(n5504) );
  DFE1 \mem_reg_26][15  ( .D(D_15), .E(n6451), .C(wclk), .QN(n5505) );
  DFE1 \mem_reg_26][14  ( .D(D_14), .E(n6451), .C(wclk), .QN(n5506) );
  DFE1 \mem_reg_26][13  ( .D(D_13), .E(n6451), .C(wclk), .QN(n5507) );
  DFE1 \mem_reg_26][12  ( .D(D_12), .E(n6451), .C(wclk), .QN(n5508) );
  DFE1 \mem_reg_26][11  ( .D(D_11), .E(n6451), .C(wclk), .QN(n5509) );
  DFE1 \mem_reg_26][10  ( .D(D_10), .E(n6451), .C(wclk), .QN(n5510) );
  DFE1 \mem_reg_26][9  ( .D(D_9), .E(n6451), .C(wclk), .QN(n5511) );
  DFE1 \mem_reg_26][8  ( .D(D_8), .E(n6451), .C(wclk), .QN(n5512) );
  DFE1 \mem_reg_26][7  ( .D(D_7), .E(n6451), .C(wclk), .QN(n5513) );
  DFE1 \mem_reg_26][6  ( .D(D_6), .E(n6451), .C(wclk), .QN(n5514) );
  DFE1 \mem_reg_26][5  ( .D(D_5), .E(n6451), .C(wclk), .QN(n5515) );
  DFE1 \mem_reg_26][4  ( .D(D_4), .E(n6451), .C(wclk), .QN(n5516) );
  DFE1 \mem_reg_26][3  ( .D(D_3), .E(n6451), .C(wclk), .QN(n5517) );
  DFE1 \mem_reg_26][2  ( .D(D_2), .E(n6451), .C(wclk), .QN(n5518) );
  DFE1 \mem_reg_26][1  ( .D(D_1), .E(n6451), .C(wclk), .QN(n5519) );
  DFE1 \mem_reg_26][0  ( .D(D_0), .E(n6451), .C(wclk), .QN(n5520) );
  DFE1 \mem_reg_25][23  ( .D(D_23), .E(n6450), .C(wclk), .QN(n5521) );
  DFE1 \mem_reg_25][22  ( .D(D_22), .E(n6450), .C(wclk), .QN(n5522) );
  DFE1 \mem_reg_25][21  ( .D(D_21), .E(n6450), .C(wclk), .QN(n5523) );
  DFE1 \mem_reg_25][20  ( .D(D_20), .E(n6450), .C(wclk), .QN(n5524) );
  DFE1 \mem_reg_25][19  ( .D(D_19), .E(n6450), .C(wclk), .QN(n5525) );
  DFE1 \mem_reg_25][18  ( .D(D_18), .E(n6450), .C(wclk), .QN(n5526) );
  DFE1 \mem_reg_25][17  ( .D(D_17), .E(n6450), .C(wclk), .QN(n5527) );
  DFE1 \mem_reg_25][16  ( .D(D_16), .E(n6450), .C(wclk), .QN(n5528) );
  DFE1 \mem_reg_25][15  ( .D(D_15), .E(n6450), .C(wclk), .QN(n5529) );
  DFE1 \mem_reg_25][14  ( .D(D_14), .E(n6450), .C(wclk), .QN(n5530) );
  DFE1 \mem_reg_25][13  ( .D(D_13), .E(n6450), .C(wclk), .QN(n5531) );
  DFE1 \mem_reg_25][12  ( .D(D_12), .E(n6450), .C(wclk), .QN(n5532) );
  DFE1 \mem_reg_25][11  ( .D(D_11), .E(n6450), .C(wclk), .QN(n5533) );
  DFE1 \mem_reg_25][10  ( .D(D_10), .E(n6450), .C(wclk), .QN(n5534) );
  DFE1 \mem_reg_25][9  ( .D(D_9), .E(n6450), .C(wclk), .QN(n5535) );
  DFE1 \mem_reg_25][8  ( .D(D_8), .E(n6450), .C(wclk), .QN(n5536) );
  DFE1 \mem_reg_25][7  ( .D(D_7), .E(n6450), .C(wclk), .QN(n5537) );
  DFE1 \mem_reg_25][6  ( .D(D_6), .E(n6450), .C(wclk), .QN(n5538) );
  DFE1 \mem_reg_25][5  ( .D(D_5), .E(n6450), .C(wclk), .QN(n5539) );
  DFE1 \mem_reg_25][4  ( .D(D_4), .E(n6450), .C(wclk), .QN(n5540) );
  DFE1 \mem_reg_25][3  ( .D(D_3), .E(n6450), .C(wclk), .QN(n5541) );
  DFE1 \mem_reg_25][2  ( .D(D_2), .E(n6450), .C(wclk), .QN(n5542) );
  DFE1 \mem_reg_25][1  ( .D(D_1), .E(n6450), .C(wclk), .QN(n5543) );
  DFE1 \mem_reg_25][0  ( .D(D_0), .E(n6450), .C(wclk), .QN(n5544) );
  DFE1 \mem_reg_24][23  ( .D(D_23), .E(n6449), .C(wclk), .QN(n5545) );
  DFE1 \mem_reg_24][22  ( .D(D_22), .E(n6449), .C(wclk), .QN(n5546) );
  DFE1 \mem_reg_24][21  ( .D(D_21), .E(n6449), .C(wclk), .QN(n5547) );
  DFE1 \mem_reg_24][20  ( .D(D_20), .E(n6449), .C(wclk), .QN(n5548) );
  DFE1 \mem_reg_24][19  ( .D(D_19), .E(n6449), .C(wclk), .QN(n5549) );
  DFE1 \mem_reg_24][18  ( .D(D_18), .E(n6449), .C(wclk), .QN(n5550) );
  DFE1 \mem_reg_24][17  ( .D(D_17), .E(n6449), .C(wclk), .QN(n5551) );
  DFE1 \mem_reg_24][16  ( .D(D_16), .E(n6449), .C(wclk), .QN(n5552) );
  DFE1 \mem_reg_24][15  ( .D(D_15), .E(n6449), .C(wclk), .QN(n5553) );
  DFE1 \mem_reg_24][14  ( .D(D_14), .E(n6449), .C(wclk), .QN(n5554) );
  DFE1 \mem_reg_24][13  ( .D(D_13), .E(n6449), .C(wclk), .QN(n5555) );
  DFE1 \mem_reg_24][12  ( .D(D_12), .E(n6449), .C(wclk), .QN(n5556) );
  DFE1 \mem_reg_24][11  ( .D(D_11), .E(n6449), .C(wclk), .QN(n5557) );
  DFE1 \mem_reg_24][10  ( .D(D_10), .E(n6449), .C(wclk), .QN(n5558) );
  DFE1 \mem_reg_24][9  ( .D(D_9), .E(n6449), .C(wclk), .QN(n5559) );
  DFE1 \mem_reg_24][8  ( .D(D_8), .E(n6449), .C(wclk), .QN(n5560) );
  DFE1 \mem_reg_24][7  ( .D(D_7), .E(n6449), .C(wclk), .QN(n5561) );
  DFE1 \mem_reg_24][6  ( .D(D_6), .E(n6449), .C(wclk), .QN(n5562) );
  DFE1 \mem_reg_24][5  ( .D(D_5), .E(n6449), .C(wclk), .QN(n5563) );
  DFE1 \mem_reg_24][4  ( .D(D_4), .E(n6449), .C(wclk), .QN(n5564) );
  DFE1 \mem_reg_24][3  ( .D(D_3), .E(n6449), .C(wclk), .QN(n5565) );
  DFE1 \mem_reg_24][2  ( .D(D_2), .E(n6449), .C(wclk), .QN(n5566) );
  DFE1 \mem_reg_24][1  ( .D(D_1), .E(n6449), .C(wclk), .QN(n5567) );
  DFE1 \mem_reg_24][0  ( .D(D_0), .E(n6449), .C(wclk), .QN(n5568) );
  DFE1 \mem_reg_23][23  ( .D(D_23), .E(n6447), .C(wclk), .QN(n5569) );
  DFE1 \mem_reg_23][22  ( .D(D_22), .E(n6447), .C(wclk), .QN(n5570) );
  DFE1 \mem_reg_23][21  ( .D(D_21), .E(n6447), .C(wclk), .QN(n5571) );
  DFE1 \mem_reg_23][20  ( .D(D_20), .E(n6447), .C(wclk), .QN(n5572) );
  DFE1 \mem_reg_23][19  ( .D(D_19), .E(n6447), .C(wclk), .QN(n5573) );
  DFE1 \mem_reg_23][18  ( .D(D_18), .E(n6447), .C(wclk), .QN(n5574) );
  DFE1 \mem_reg_23][17  ( .D(D_17), .E(n6447), .C(wclk), .QN(n5575) );
  DFE1 \mem_reg_23][16  ( .D(D_16), .E(n6447), .C(wclk), .QN(n5576) );
  DFE1 \mem_reg_23][15  ( .D(D_15), .E(n6447), .C(wclk), .QN(n5577) );
  DFE1 \mem_reg_23][14  ( .D(D_14), .E(n6447), .C(wclk), .QN(n5578) );
  DFE1 \mem_reg_23][13  ( .D(D_13), .E(n6447), .C(wclk), .QN(n5579) );
  DFE1 \mem_reg_23][12  ( .D(D_12), .E(n6447), .C(wclk), .QN(n5580) );
  DFE1 \mem_reg_23][11  ( .D(D_11), .E(n6447), .C(wclk), .QN(n5581) );
  DFE1 \mem_reg_23][10  ( .D(D_10), .E(n6447), .C(wclk), .QN(n5582) );
  DFE1 \mem_reg_23][9  ( .D(D_9), .E(n6447), .C(wclk), .QN(n5583) );
  DFE1 \mem_reg_23][8  ( .D(D_8), .E(n6447), .C(wclk), .QN(n5584) );
  DFE1 \mem_reg_23][7  ( .D(D_7), .E(n6447), .C(wclk), .QN(n5585) );
  DFE1 \mem_reg_23][6  ( .D(D_6), .E(n6447), .C(wclk), .QN(n5586) );
  DFE1 \mem_reg_23][5  ( .D(D_5), .E(n6447), .C(wclk), .QN(n5587) );
  DFE1 \mem_reg_23][4  ( .D(D_4), .E(n6447), .C(wclk), .QN(n5588) );
  DFE1 \mem_reg_23][3  ( .D(D_3), .E(n6447), .C(wclk), .QN(n5589) );
  DFE1 \mem_reg_23][2  ( .D(D_2), .E(n6447), .C(wclk), .QN(n5590) );
  DFE1 \mem_reg_23][1  ( .D(D_1), .E(n6447), .C(wclk), .QN(n5591) );
  DFE1 \mem_reg_23][0  ( .D(D_0), .E(n6447), .C(wclk), .QN(n5592) );
  DFE1 \mem_reg_22][23  ( .D(D_23), .E(n6446), .C(wclk), .QN(n5593) );
  DFE1 \mem_reg_22][22  ( .D(D_22), .E(n6446), .C(wclk), .QN(n5594) );
  DFE1 \mem_reg_22][21  ( .D(D_21), .E(n6446), .C(wclk), .QN(n5595) );
  DFE1 \mem_reg_22][20  ( .D(D_20), .E(n6446), .C(wclk), .QN(n5596) );
  DFE1 \mem_reg_22][19  ( .D(D_19), .E(n6446), .C(wclk), .QN(n5597) );
  DFE1 \mem_reg_22][18  ( .D(D_18), .E(n6446), .C(wclk), .QN(n5598) );
  DFE1 \mem_reg_22][17  ( .D(D_17), .E(n6446), .C(wclk), .QN(n5599) );
  DFE1 \mem_reg_22][16  ( .D(D_16), .E(n6446), .C(wclk), .QN(n5600) );
  DFE1 \mem_reg_22][15  ( .D(D_15), .E(n6446), .C(wclk), .QN(n5601) );
  DFE1 \mem_reg_22][14  ( .D(D_14), .E(n6446), .C(wclk), .QN(n5602) );
  DFE1 \mem_reg_22][13  ( .D(D_13), .E(n6446), .C(wclk), .QN(n5603) );
  DFE1 \mem_reg_22][12  ( .D(D_12), .E(n6446), .C(wclk), .QN(n5604) );
  DFE1 \mem_reg_22][11  ( .D(D_11), .E(n6446), .C(wclk), .QN(n5605) );
  DFE1 \mem_reg_22][10  ( .D(D_10), .E(n6446), .C(wclk), .QN(n5606) );
  DFE1 \mem_reg_22][9  ( .D(D_9), .E(n6446), .C(wclk), .QN(n5607) );
  DFE1 \mem_reg_22][8  ( .D(D_8), .E(n6446), .C(wclk), .QN(n5608) );
  DFE1 \mem_reg_22][7  ( .D(D_7), .E(n6446), .C(wclk), .QN(n5609) );
  DFE1 \mem_reg_22][6  ( .D(D_6), .E(n6446), .C(wclk), .QN(n5610) );
  DFE1 \mem_reg_22][5  ( .D(D_5), .E(n6446), .C(wclk), .QN(n5611) );
  DFE1 \mem_reg_22][4  ( .D(D_4), .E(n6446), .C(wclk), .QN(n5612) );
  DFE1 \mem_reg_22][3  ( .D(D_3), .E(n6446), .C(wclk), .QN(n5613) );
  DFE1 \mem_reg_22][2  ( .D(D_2), .E(n6446), .C(wclk), .QN(n5614) );
  DFE1 \mem_reg_22][1  ( .D(D_1), .E(n6446), .C(wclk), .QN(n5615) );
  DFE1 \mem_reg_22][0  ( .D(D_0), .E(n6446), .C(wclk), .QN(n5616) );
  DFE1 \mem_reg_21][23  ( .D(D_23), .E(n6445), .C(wclk), .QN(n5617) );
  DFE1 \mem_reg_21][22  ( .D(D_22), .E(n6445), .C(wclk), .QN(n5618) );
  DFE1 \mem_reg_21][21  ( .D(D_21), .E(n6445), .C(wclk), .QN(n5619) );
  DFE1 \mem_reg_21][20  ( .D(D_20), .E(n6445), .C(wclk), .QN(n5620) );
  DFE1 \mem_reg_21][19  ( .D(D_19), .E(n6445), .C(wclk), .QN(n5621) );
  DFE1 \mem_reg_21][18  ( .D(D_18), .E(n6445), .C(wclk), .QN(n5622) );
  DFE1 \mem_reg_21][17  ( .D(D_17), .E(n6445), .C(wclk), .QN(n5623) );
  DFE1 \mem_reg_21][16  ( .D(D_16), .E(n6445), .C(wclk), .QN(n5624) );
  DFE1 \mem_reg_21][15  ( .D(D_15), .E(n6445), .C(wclk), .QN(n5625) );
  DFE1 \mem_reg_21][14  ( .D(D_14), .E(n6445), .C(wclk), .QN(n5626) );
  DFE1 \mem_reg_21][13  ( .D(D_13), .E(n6445), .C(wclk), .QN(n5627) );
  DFE1 \mem_reg_21][12  ( .D(D_12), .E(n6445), .C(wclk), .QN(n5628) );
  DFE1 \mem_reg_21][11  ( .D(D_11), .E(n6445), .C(wclk), .QN(n5629) );
  DFE1 \mem_reg_21][10  ( .D(D_10), .E(n6445), .C(wclk), .QN(n5630) );
  DFE1 \mem_reg_21][9  ( .D(D_9), .E(n6445), .C(wclk), .QN(n5631) );
  DFE1 \mem_reg_21][8  ( .D(D_8), .E(n6445), .C(wclk), .QN(n5632) );
  DFE1 \mem_reg_21][7  ( .D(D_7), .E(n6445), .C(wclk), .QN(n5633) );
  DFE1 \mem_reg_21][6  ( .D(D_6), .E(n6445), .C(wclk), .QN(n5634) );
  DFE1 \mem_reg_21][5  ( .D(D_5), .E(n6445), .C(wclk), .QN(n5635) );
  DFE1 \mem_reg_21][4  ( .D(D_4), .E(n6445), .C(wclk), .QN(n5636) );
  DFE1 \mem_reg_21][3  ( .D(D_3), .E(n6445), .C(wclk), .QN(n5637) );
  DFE1 \mem_reg_21][2  ( .D(D_2), .E(n6445), .C(wclk), .QN(n5638) );
  DFE1 \mem_reg_21][1  ( .D(D_1), .E(n6445), .C(wclk), .QN(n5639) );
  DFE1 \mem_reg_21][0  ( .D(D_0), .E(n6445), .C(wclk), .QN(n5640) );
  DFE1 \mem_reg_20][23  ( .D(D_23), .E(n6444), .C(wclk), .QN(n5641) );
  DFE1 \mem_reg_20][22  ( .D(D_22), .E(n6444), .C(wclk), .QN(n5642) );
  DFE1 \mem_reg_20][21  ( .D(D_21), .E(n6444), .C(wclk), .QN(n5643) );
  DFE1 \mem_reg_20][20  ( .D(D_20), .E(n6444), .C(wclk), .QN(n5644) );
  DFE1 \mem_reg_20][19  ( .D(D_19), .E(n6444), .C(wclk), .QN(n5645) );
  DFE1 \mem_reg_20][18  ( .D(D_18), .E(n6444), .C(wclk), .QN(n5646) );
  DFE1 \mem_reg_20][17  ( .D(D_17), .E(n6444), .C(wclk), .QN(n5647) );
  DFE1 \mem_reg_20][16  ( .D(D_16), .E(n6444), .C(wclk), .QN(n5648) );
  DFE1 \mem_reg_20][15  ( .D(D_15), .E(n6444), .C(wclk), .QN(n5649) );
  DFE1 \mem_reg_20][14  ( .D(D_14), .E(n6444), .C(wclk), .QN(n5650) );
  DFE1 \mem_reg_20][13  ( .D(D_13), .E(n6444), .C(wclk), .QN(n5651) );
  DFE1 \mem_reg_20][12  ( .D(D_12), .E(n6444), .C(wclk), .QN(n5652) );
  DFE1 \mem_reg_20][11  ( .D(D_11), .E(n6444), .C(wclk), .QN(n5653) );
  DFE1 \mem_reg_20][10  ( .D(D_10), .E(n6444), .C(wclk), .QN(n5654) );
  DFE1 \mem_reg_20][9  ( .D(D_9), .E(n6444), .C(wclk), .QN(n5655) );
  DFE1 \mem_reg_20][8  ( .D(D_8), .E(n6444), .C(wclk), .QN(n5656) );
  DFE1 \mem_reg_20][7  ( .D(D_7), .E(n6444), .C(wclk), .QN(n5657) );
  DFE1 \mem_reg_20][6  ( .D(D_6), .E(n6444), .C(wclk), .QN(n5658) );
  DFE1 \mem_reg_20][5  ( .D(D_5), .E(n6444), .C(wclk), .QN(n5659) );
  DFE1 \mem_reg_20][4  ( .D(D_4), .E(n6444), .C(wclk), .QN(n5660) );
  DFE1 \mem_reg_20][3  ( .D(D_3), .E(n6444), .C(wclk), .QN(n5661) );
  DFE1 \mem_reg_20][2  ( .D(D_2), .E(n6444), .C(wclk), .QN(n5662) );
  DFE1 \mem_reg_20][1  ( .D(D_1), .E(n6444), .C(wclk), .QN(n5663) );
  DFE1 \mem_reg_20][0  ( .D(D_0), .E(n6444), .C(wclk), .QN(n5664) );
  DFE1 \mem_reg_19][23  ( .D(D_23), .E(n6443), .C(wclk), .QN(n5665) );
  DFE1 \mem_reg_19][22  ( .D(D_22), .E(n6443), .C(wclk), .QN(n5666) );
  DFE1 \mem_reg_19][21  ( .D(D_21), .E(n6443), .C(wclk), .QN(n5667) );
  DFE1 \mem_reg_19][20  ( .D(D_20), .E(n6443), .C(wclk), .QN(n5668) );
  DFE1 \mem_reg_19][19  ( .D(D_19), .E(n6443), .C(wclk), .QN(n5669) );
  DFE1 \mem_reg_19][18  ( .D(D_18), .E(n6443), .C(wclk), .QN(n5670) );
  DFE1 \mem_reg_19][17  ( .D(D_17), .E(n6443), .C(wclk), .QN(n5671) );
  DFE1 \mem_reg_19][16  ( .D(D_16), .E(n6443), .C(wclk), .QN(n5672) );
  DFE1 \mem_reg_19][15  ( .D(D_15), .E(n6443), .C(wclk), .QN(n5673) );
  DFE1 \mem_reg_19][14  ( .D(D_14), .E(n6443), .C(wclk), .QN(n5674) );
  DFE1 \mem_reg_19][13  ( .D(D_13), .E(n6443), .C(wclk), .QN(n5675) );
  DFE1 \mem_reg_19][12  ( .D(D_12), .E(n6443), .C(wclk), .QN(n5676) );
  DFE1 \mem_reg_19][11  ( .D(D_11), .E(n6443), .C(wclk), .QN(n5677) );
  DFE1 \mem_reg_19][10  ( .D(D_10), .E(n6443), .C(wclk), .QN(n5678) );
  DFE1 \mem_reg_19][9  ( .D(D_9), .E(n6443), .C(wclk), .QN(n5679) );
  DFE1 \mem_reg_19][8  ( .D(D_8), .E(n6443), .C(wclk), .QN(n5680) );
  DFE1 \mem_reg_19][7  ( .D(D_7), .E(n6443), .C(wclk), .QN(n5681) );
  DFE1 \mem_reg_19][6  ( .D(D_6), .E(n6443), .C(wclk), .QN(n5682) );
  DFE1 \mem_reg_19][5  ( .D(D_5), .E(n6443), .C(wclk), .QN(n5683) );
  DFE1 \mem_reg_19][4  ( .D(D_4), .E(n6443), .C(wclk), .QN(n5684) );
  DFE1 \mem_reg_19][3  ( .D(D_3), .E(n6443), .C(wclk), .QN(n5685) );
  DFE1 \mem_reg_19][2  ( .D(D_2), .E(n6443), .C(wclk), .QN(n5686) );
  DFE1 \mem_reg_19][1  ( .D(D_1), .E(n6443), .C(wclk), .QN(n5687) );
  DFE1 \mem_reg_19][0  ( .D(D_0), .E(n6443), .C(wclk), .QN(n5688) );
  DFE1 \mem_reg_18][23  ( .D(D_23), .E(n6442), .C(wclk), .QN(n5689) );
  DFE1 \mem_reg_18][22  ( .D(D_22), .E(n6442), .C(wclk), .QN(n5690) );
  DFE1 \mem_reg_18][21  ( .D(D_21), .E(n6442), .C(wclk), .QN(n5691) );
  DFE1 \mem_reg_18][20  ( .D(D_20), .E(n6442), .C(wclk), .QN(n5692) );
  DFE1 \mem_reg_18][19  ( .D(D_19), .E(n6442), .C(wclk), .QN(n5693) );
  DFE1 \mem_reg_18][18  ( .D(D_18), .E(n6442), .C(wclk), .QN(n5694) );
  DFE1 \mem_reg_18][17  ( .D(D_17), .E(n6442), .C(wclk), .QN(n5695) );
  DFE1 \mem_reg_18][16  ( .D(D_16), .E(n6442), .C(wclk), .QN(n5696) );
  DFE1 \mem_reg_18][15  ( .D(D_15), .E(n6442), .C(wclk), .QN(n5697) );
  DFE1 \mem_reg_18][14  ( .D(D_14), .E(n6442), .C(wclk), .QN(n5698) );
  DFE1 \mem_reg_18][13  ( .D(D_13), .E(n6442), .C(wclk), .QN(n5699) );
  DFE1 \mem_reg_18][12  ( .D(D_12), .E(n6442), .C(wclk), .QN(n5700) );
  DFE1 \mem_reg_18][11  ( .D(D_11), .E(n6442), .C(wclk), .QN(n5701) );
  DFE1 \mem_reg_18][10  ( .D(D_10), .E(n6442), .C(wclk), .QN(n5702) );
  DFE1 \mem_reg_18][9  ( .D(D_9), .E(n6442), .C(wclk), .QN(n5703) );
  DFE1 \mem_reg_18][8  ( .D(D_8), .E(n6442), .C(wclk), .QN(n5704) );
  DFE1 \mem_reg_18][7  ( .D(D_7), .E(n6442), .C(wclk), .QN(n5705) );
  DFE1 \mem_reg_18][6  ( .D(D_6), .E(n6442), .C(wclk), .QN(n5706) );
  DFE1 \mem_reg_18][5  ( .D(D_5), .E(n6442), .C(wclk), .QN(n5707) );
  DFE1 \mem_reg_18][4  ( .D(D_4), .E(n6442), .C(wclk), .QN(n5708) );
  DFE1 \mem_reg_18][3  ( .D(D_3), .E(n6442), .C(wclk), .QN(n5709) );
  DFE1 \mem_reg_18][2  ( .D(D_2), .E(n6442), .C(wclk), .QN(n5710) );
  DFE1 \mem_reg_18][1  ( .D(D_1), .E(n6442), .C(wclk), .QN(n5711) );
  DFE1 \mem_reg_18][0  ( .D(D_0), .E(n6442), .C(wclk), .QN(n5712) );
  DFE1 \mem_reg_17][23  ( .D(D_23), .E(n6441), .C(wclk), .QN(n5713) );
  DFE1 \mem_reg_17][22  ( .D(D_22), .E(n6441), .C(wclk), .QN(n5714) );
  DFE1 \mem_reg_17][21  ( .D(D_21), .E(n6441), .C(wclk), .QN(n5715) );
  DFE1 \mem_reg_17][20  ( .D(D_20), .E(n6441), .C(wclk), .QN(n5716) );
  DFE1 \mem_reg_17][19  ( .D(D_19), .E(n6441), .C(wclk), .QN(n5717) );
  DFE1 \mem_reg_17][18  ( .D(D_18), .E(n6441), .C(wclk), .QN(n5718) );
  DFE1 \mem_reg_17][17  ( .D(D_17), .E(n6441), .C(wclk), .QN(n5719) );
  DFE1 \mem_reg_17][16  ( .D(D_16), .E(n6441), .C(wclk), .QN(n5720) );
  DFE1 \mem_reg_17][15  ( .D(D_15), .E(n6441), .C(wclk), .QN(n5721) );
  DFE1 \mem_reg_17][14  ( .D(D_14), .E(n6441), .C(wclk), .QN(n5722) );
  DFE1 \mem_reg_17][13  ( .D(D_13), .E(n6441), .C(wclk), .QN(n5723) );
  DFE1 \mem_reg_17][12  ( .D(D_12), .E(n6441), .C(wclk), .QN(n5724) );
  DFE1 \mem_reg_17][11  ( .D(D_11), .E(n6441), .C(wclk), .QN(n5725) );
  DFE1 \mem_reg_17][10  ( .D(D_10), .E(n6441), .C(wclk), .QN(n5726) );
  DFE1 \mem_reg_17][9  ( .D(D_9), .E(n6441), .C(wclk), .QN(n5727) );
  DFE1 \mem_reg_17][8  ( .D(D_8), .E(n6441), .C(wclk), .QN(n5728) );
  DFE1 \mem_reg_17][7  ( .D(D_7), .E(n6441), .C(wclk), .QN(n5729) );
  DFE1 \mem_reg_17][6  ( .D(D_6), .E(n6441), .C(wclk), .QN(n5730) );
  DFE1 \mem_reg_17][5  ( .D(D_5), .E(n6441), .C(wclk), .QN(n5731) );
  DFE1 \mem_reg_17][4  ( .D(D_4), .E(n6441), .C(wclk), .QN(n5732) );
  DFE1 \mem_reg_17][3  ( .D(D_3), .E(n6441), .C(wclk), .QN(n5733) );
  DFE1 \mem_reg_17][2  ( .D(D_2), .E(n6441), .C(wclk), .QN(n5734) );
  DFE1 \mem_reg_17][1  ( .D(D_1), .E(n6441), .C(wclk), .QN(n5735) );
  DFE1 \mem_reg_17][0  ( .D(D_0), .E(n6441), .C(wclk), .QN(n5736) );
  DFE1 \mem_reg_16][23  ( .D(D_23), .E(n6439), .C(wclk), .QN(n5737) );
  DFE1 \mem_reg_16][22  ( .D(D_22), .E(n6439), .C(wclk), .QN(n5738) );
  DFE1 \mem_reg_16][21  ( .D(D_21), .E(n6439), .C(wclk), .QN(n5739) );
  DFE1 \mem_reg_16][20  ( .D(D_20), .E(n6439), .C(wclk), .QN(n5740) );
  DFE1 \mem_reg_16][19  ( .D(D_19), .E(n6439), .C(wclk), .QN(n5741) );
  DFE1 \mem_reg_16][18  ( .D(D_18), .E(n6439), .C(wclk), .QN(n5742) );
  DFE1 \mem_reg_16][17  ( .D(D_17), .E(n6439), .C(wclk), .QN(n5743) );
  DFE1 \mem_reg_16][16  ( .D(D_16), .E(n6439), .C(wclk), .QN(n5744) );
  DFE1 \mem_reg_16][15  ( .D(D_15), .E(n6439), .C(wclk), .QN(n5745) );
  DFE1 \mem_reg_16][14  ( .D(D_14), .E(n6439), .C(wclk), .QN(n5746) );
  DFE1 \mem_reg_16][13  ( .D(D_13), .E(n6439), .C(wclk), .QN(n5747) );
  DFE1 \mem_reg_16][12  ( .D(D_12), .E(n6439), .C(wclk), .QN(n5748) );
  DFE1 \mem_reg_16][11  ( .D(D_11), .E(n6439), .C(wclk), .QN(n5749) );
  DFE1 \mem_reg_16][10  ( .D(D_10), .E(n6439), .C(wclk), .QN(n5750) );
  DFE1 \mem_reg_16][9  ( .D(D_9), .E(n6439), .C(wclk), .QN(n5751) );
  DFE1 \mem_reg_16][8  ( .D(D_8), .E(n6439), .C(wclk), .QN(n5752) );
  DFE1 \mem_reg_16][7  ( .D(D_7), .E(n6439), .C(wclk), .QN(n5753) );
  DFE1 \mem_reg_16][6  ( .D(D_6), .E(n6439), .C(wclk), .QN(n5754) );
  DFE1 \mem_reg_16][5  ( .D(D_5), .E(n6439), .C(wclk), .QN(n5755) );
  DFE1 \mem_reg_16][4  ( .D(D_4), .E(n6439), .C(wclk), .QN(n5756) );
  DFE1 \mem_reg_16][3  ( .D(D_3), .E(n6439), .C(wclk), .QN(n5757) );
  DFE1 \mem_reg_16][2  ( .D(D_2), .E(n6439), .C(wclk), .QN(n5758) );
  DFE1 \mem_reg_16][1  ( .D(D_1), .E(n6439), .C(wclk), .QN(n5759) );
  DFE1 \mem_reg_16][0  ( .D(D_0), .E(n6439), .C(wclk), .QN(n5760) );
  NOR21 U3 ( .A(waddr_5), .B(waddr_4), .Q(n6234) );
  NOR23 U4 ( .A(n11159), .B(n11135), .Q(n6313) );
  NOR23 U5 ( .A(n11159), .B(n11131), .Q(n6315) );
  NOR23 U6 ( .A(n11159), .B(n11128), .Q(n6316) );
  NOR23 U7 ( .A(n11159), .B(n11125), .Q(n6317) );
  NOR23 U8 ( .A(n11159), .B(n11122), .Q(n6318) );
  NOR23 U9 ( .A(n11159), .B(n11119), .Q(n6319) );
  NOR23 U10 ( .A(n11159), .B(n11116), .Q(n6320) );
  NOR23 U11 ( .A(n11159), .B(n11113), .Q(n6321) );
  CLKBU2 U12 ( .A(n6314), .Q(n11159) );
  NOR23 U13 ( .A(n11158), .B(n11101), .Q(n6322) );
  NOR23 U14 ( .A(n11158), .B(n11111), .Q(n6323) );
  NOR23 U15 ( .A(n11158), .B(n11108), .Q(n6324) );
  NOR23 U16 ( .A(n11158), .B(n11106), .Q(n6325) );
  NOR23 U17 ( .A(n11158), .B(n11103), .Q(n6326) );
  NOR23 U18 ( .A(n11158), .B(n11095), .Q(n6327) );
  NOR23 U19 ( .A(n11158), .B(n11143), .Q(n6328) );
  NOR23 U20 ( .A(n11158), .B(n11140), .Q(n6329) );
  CLKBU2 U21 ( .A(n6314), .Q(n11158) );
  NOR23 U22 ( .A(n11157), .B(n11134), .Q(n6330) );
  NOR23 U23 ( .A(n11157), .B(n11132), .Q(n6332) );
  NOR23 U24 ( .A(n11157), .B(n11129), .Q(n6333) );
  NOR23 U25 ( .A(n11157), .B(n11126), .Q(n6334) );
  NOR23 U26 ( .A(n11157), .B(n11123), .Q(n6335) );
  NOR23 U27 ( .A(n11157), .B(n11120), .Q(n6336) );
  NOR23 U28 ( .A(n11157), .B(n11117), .Q(n6337) );
  NOR23 U29 ( .A(n11157), .B(n11114), .Q(n6338) );
  CLKBU2 U30 ( .A(n6331), .Q(n11157) );
  NOR23 U31 ( .A(n11156), .B(n11100), .Q(n6339) );
  NOR23 U32 ( .A(n11156), .B(n11110), .Q(n6340) );
  NOR23 U33 ( .A(n11156), .B(n11108), .Q(n6341) );
  NOR23 U34 ( .A(n11156), .B(n11106), .Q(n6342) );
  NOR23 U35 ( .A(n11156), .B(n11104), .Q(n6343) );
  NOR23 U36 ( .A(n11156), .B(n11096), .Q(n6344) );
  NOR23 U37 ( .A(n11156), .B(n11142), .Q(n6345) );
  NOR23 U38 ( .A(n11156), .B(n11139), .Q(n6346) );
  CLKBU2 U39 ( .A(n6331), .Q(n11156) );
  NOR23 U40 ( .A(n11167), .B(n11135), .Q(n6236) );
  NOR23 U41 ( .A(n11167), .B(n11131), .Q(n6238) );
  NOR23 U42 ( .A(n11167), .B(n11128), .Q(n6239) );
  NOR23 U43 ( .A(n11167), .B(n11125), .Q(n6240) );
  NOR23 U44 ( .A(n11167), .B(n11122), .Q(n6242) );
  NOR23 U45 ( .A(n11167), .B(n11119), .Q(n6243) );
  CLKBU2 U46 ( .A(n6213), .Q(n11119) );
  NOR23 U47 ( .A(n11167), .B(n11116), .Q(n6244) );
  NOR23 U48 ( .A(n11167), .B(n11113), .Q(n6245) );
  CLKBU2 U49 ( .A(n6237), .Q(n11167) );
  NOR23 U50 ( .A(n11166), .B(n11101), .Q(n6246) );
  NOR23 U51 ( .A(n11166), .B(n11111), .Q(n6247) );
  NOR23 U52 ( .A(n11166), .B(n11108), .Q(n6248) );
  NOR23 U53 ( .A(n11166), .B(n11106), .Q(n6249) );
  NOR23 U54 ( .A(n11166), .B(n11103), .Q(n6250) );
  NOR23 U55 ( .A(n11166), .B(n11096), .Q(n6251) );
  NOR23 U56 ( .A(n11166), .B(n11143), .Q(n6253) );
  NOR23 U57 ( .A(n11166), .B(n11140), .Q(n6254) );
  CLKBU2 U58 ( .A(n6237), .Q(n11166) );
  NOR23 U59 ( .A(n11165), .B(n11134), .Q(n6256) );
  NOR23 U60 ( .A(n11165), .B(n11132), .Q(n6258) );
  NOR23 U61 ( .A(n11165), .B(n11129), .Q(n6259) );
  NOR23 U62 ( .A(n11165), .B(n11126), .Q(n6260) );
  NOR23 U63 ( .A(n11165), .B(n11123), .Q(n6261) );
  NOR23 U64 ( .A(n11165), .B(n11120), .Q(n6262) );
  NOR23 U65 ( .A(n11165), .B(n11117), .Q(n6263) );
  NOR23 U66 ( .A(n11165), .B(n11114), .Q(n6264) );
  CLKBU2 U67 ( .A(n6257), .Q(n11165) );
  NOR23 U68 ( .A(n11164), .B(n11100), .Q(n6266) );
  NOR23 U69 ( .A(n11164), .B(n11110), .Q(n6267) );
  NOR23 U70 ( .A(n11164), .B(n11108), .Q(n6268) );
  NOR23 U71 ( .A(n11164), .B(n11106), .Q(n6269) );
  NOR23 U72 ( .A(n11164), .B(n11104), .Q(n6270) );
  NOR23 U73 ( .A(n11164), .B(n11095), .Q(n6271) );
  NOR23 U74 ( .A(n11164), .B(n11142), .Q(n6272) );
  NOR23 U75 ( .A(n11164), .B(n11139), .Q(n6273) );
  CLKBU2 U76 ( .A(n6257), .Q(n11164) );
  NOR23 U77 ( .A(n11161), .B(n11134), .Q(n6295) );
  NOR23 U78 ( .A(n11161), .B(n11132), .Q(n6297) );
  NOR23 U79 ( .A(n11161), .B(n11129), .Q(n6298) );
  NOR23 U80 ( .A(n11161), .B(n11126), .Q(n6299) );
  NOR23 U81 ( .A(n11161), .B(n11123), .Q(n6300) );
  NOR23 U82 ( .A(n11161), .B(n11120), .Q(n6301) );
  NOR23 U83 ( .A(n11161), .B(n11117), .Q(n6302) );
  CLKBU2 U84 ( .A(n6215), .Q(n11117) );
  NOR23 U85 ( .A(n11161), .B(n11114), .Q(n6303) );
  CLKBU2 U86 ( .A(n6296), .Q(n11161) );
  NOR23 U87 ( .A(n11160), .B(n11100), .Q(n6304) );
  NOR23 U88 ( .A(n11160), .B(n11110), .Q(n6305) );
  NOR23 U89 ( .A(n11160), .B(n11108), .Q(n6306) );
  CLKBU2 U90 ( .A(n6225), .Q(n11108) );
  NOR23 U91 ( .A(n11160), .B(n11106), .Q(n6307) );
  CLKBU2 U92 ( .A(n6227), .Q(n11106) );
  NOR23 U93 ( .A(n11160), .B(n11104), .Q(n6308) );
  NOR23 U94 ( .A(n11160), .B(n11096), .Q(n6309) );
  NOR23 U95 ( .A(n11160), .B(n11142), .Q(n6310) );
  NOR23 U96 ( .A(n11160), .B(n11139), .Q(n6311) );
  CLKBU2 U97 ( .A(n6296), .Q(n11160) );
  NOR23 U98 ( .A(n11155), .B(n11135), .Q(n6347) );
  NOR23 U99 ( .A(n11155), .B(n11131), .Q(n6349) );
  NOR23 U100 ( .A(n11155), .B(n11128), .Q(n6350) );
  NOR23 U101 ( .A(n11155), .B(n11125), .Q(n6351) );
  NOR23 U102 ( .A(n11155), .B(n11122), .Q(n6352) );
  NOR23 U103 ( .A(n11155), .B(n11119), .Q(n6353) );
  NOR23 U104 ( .A(n11155), .B(n11116), .Q(n6354) );
  NOR23 U105 ( .A(n11155), .B(n11113), .Q(n6355) );
  CLKBU2 U106 ( .A(n6348), .Q(n11155) );
  NOR23 U107 ( .A(n11154), .B(n11101), .Q(n6356) );
  NOR23 U108 ( .A(n11154), .B(n11111), .Q(n6357) );
  NOR23 U109 ( .A(n11154), .B(n11108), .Q(n6358) );
  NOR23 U110 ( .A(n11154), .B(n11106), .Q(n6359) );
  NOR23 U111 ( .A(n11154), .B(n11103), .Q(n6360) );
  NOR23 U112 ( .A(n11154), .B(n11095), .Q(n6361) );
  NOR23 U113 ( .A(n11154), .B(n11143), .Q(n6362) );
  NOR23 U114 ( .A(n11154), .B(n11140), .Q(n6363) );
  CLKBU2 U115 ( .A(n6348), .Q(n11154) );
  NOR23 U116 ( .A(n11153), .B(n11134), .Q(n6364) );
  NOR23 U117 ( .A(n11153), .B(n11132), .Q(n6366) );
  NOR23 U118 ( .A(n11153), .B(n11129), .Q(n6367) );
  NOR23 U119 ( .A(n11153), .B(n11126), .Q(n6368) );
  NOR23 U120 ( .A(n11153), .B(n11123), .Q(n6369) );
  NOR23 U121 ( .A(n11153), .B(n11120), .Q(n6370) );
  NOR23 U122 ( .A(n11153), .B(n11117), .Q(n6371) );
  NOR23 U123 ( .A(n11153), .B(n11114), .Q(n6372) );
  CLKBU2 U124 ( .A(n6217), .Q(n11114) );
  NOR23 U125 ( .A(n11152), .B(n11100), .Q(n6373) );
  NOR23 U126 ( .A(n11152), .B(n11110), .Q(n6374) );
  NOR23 U127 ( .A(n11152), .B(n11108), .Q(n6375) );
  NOR23 U128 ( .A(n11152), .B(n11106), .Q(n6376) );
  NOR23 U129 ( .A(n11152), .B(n11104), .Q(n6377) );
  NOR23 U130 ( .A(n11152), .B(n11096), .Q(n6378) );
  NOR23 U131 ( .A(n11152), .B(n11142), .Q(n6379) );
  CLKBU2 U132 ( .A(n6196), .Q(n11142) );
  NOR23 U133 ( .A(n11152), .B(n11139), .Q(n6380) );
  CLKBU2 U134 ( .A(n6365), .Q(n11152) );
  NOR23 U135 ( .A(n11151), .B(n11135), .Q(n6382) );
  NOR23 U136 ( .A(n11151), .B(n11131), .Q(n6384) );
  NOR23 U137 ( .A(n11151), .B(n11128), .Q(n6385) );
  NOR23 U138 ( .A(n11151), .B(n11125), .Q(n6386) );
  NOR23 U139 ( .A(n11151), .B(n11122), .Q(n6387) );
  NOR23 U140 ( .A(n11151), .B(n11119), .Q(n6388) );
  NOR23 U141 ( .A(n11151), .B(n11116), .Q(n6389) );
  NOR23 U142 ( .A(n11151), .B(n11113), .Q(n6390) );
  CLKBU2 U143 ( .A(n6383), .Q(n11151) );
  NOR23 U144 ( .A(n11150), .B(n11101), .Q(n6391) );
  NOR23 U145 ( .A(n11150), .B(n11111), .Q(n6392) );
  NOR23 U146 ( .A(n11150), .B(n11107), .Q(n6393) );
  NOR23 U147 ( .A(n11150), .B(n11105), .Q(n6394) );
  NOR23 U148 ( .A(n11150), .B(n11103), .Q(n6395) );
  NOR23 U149 ( .A(n11150), .B(n11094), .Q(n6396) );
  NOR23 U150 ( .A(n11150), .B(n11143), .Q(n6397) );
  NOR23 U151 ( .A(n11150), .B(n11140), .Q(n6398) );
  CLKBU2 U152 ( .A(n6383), .Q(n11150) );
  NOR23 U153 ( .A(n11149), .B(n11134), .Q(n6399) );
  NOR23 U154 ( .A(n11149), .B(n11132), .Q(n6401) );
  NOR23 U155 ( .A(n11149), .B(n11129), .Q(n6402) );
  NOR23 U156 ( .A(n11149), .B(n11126), .Q(n6403) );
  NOR23 U157 ( .A(n11149), .B(n11123), .Q(n6404) );
  NOR23 U158 ( .A(n11149), .B(n11120), .Q(n6405) );
  NOR23 U159 ( .A(n11149), .B(n11117), .Q(n6406) );
  NOR23 U160 ( .A(n11149), .B(n11114), .Q(n6407) );
  NOR23 U161 ( .A(n11148), .B(n11100), .Q(n6408) );
  NOR23 U162 ( .A(n11148), .B(n11110), .Q(n6409) );
  NOR23 U163 ( .A(n11148), .B(n11107), .Q(n6410) );
  NOR23 U164 ( .A(n11148), .B(n11105), .Q(n6411) );
  NOR23 U165 ( .A(n11148), .B(n11104), .Q(n6412) );
  NOR23 U166 ( .A(n11148), .B(n11094), .Q(n6413) );
  NOR23 U167 ( .A(n11148), .B(n11142), .Q(n6414) );
  NOR23 U168 ( .A(n11148), .B(n11139), .Q(n6415) );
  CLKBU2 U169 ( .A(n6400), .Q(n11148) );
  NOR23 U170 ( .A(n11147), .B(n11133), .Q(n6419) );
  NOR23 U171 ( .A(n11147), .B(n11131), .Q(n6421) );
  NOR23 U172 ( .A(n11147), .B(n11128), .Q(n6422) );
  NOR23 U173 ( .A(n11147), .B(n11125), .Q(n6423) );
  NOR23 U174 ( .A(n11147), .B(n11122), .Q(n6425) );
  NOR23 U175 ( .A(n11147), .B(n11119), .Q(n6426) );
  NOR23 U176 ( .A(n11147), .B(n11116), .Q(n6427) );
  NOR23 U177 ( .A(n11147), .B(n11113), .Q(n6428) );
  CLKBU2 U178 ( .A(n6420), .Q(n11147) );
  NOR23 U179 ( .A(n11146), .B(n11099), .Q(n6429) );
  NOR23 U180 ( .A(n11146), .B(n11109), .Q(n6430) );
  NOR23 U181 ( .A(n11146), .B(n11107), .Q(n6431) );
  NOR23 U182 ( .A(n11146), .B(n11105), .Q(n6432) );
  NOR23 U183 ( .A(n11146), .B(n11103), .Q(n6433) );
  NOR23 U184 ( .A(n11146), .B(n11094), .Q(n6434) );
  CLKBU2 U185 ( .A(n6231), .Q(n11094) );
  NOR23 U186 ( .A(n11146), .B(n11141), .Q(n6436) );
  NOR23 U187 ( .A(n11146), .B(n11138), .Q(n6437) );
  CLKBU2 U188 ( .A(n6420), .Q(n11146) );
  NOR23 U189 ( .A(n11145), .B(n11133), .Q(n6439) );
  NOR23 U190 ( .A(n11145), .B(n11130), .Q(n6441) );
  NOR23 U191 ( .A(n11145), .B(n11127), .Q(n6442) );
  NOR23 U192 ( .A(n11145), .B(n11124), .Q(n6443) );
  NOR23 U193 ( .A(n11145), .B(n11121), .Q(n6444) );
  NOR23 U194 ( .A(n11145), .B(n11118), .Q(n6445) );
  NOR23 U195 ( .A(n11145), .B(n11115), .Q(n6446) );
  NOR23 U196 ( .A(n11145), .B(n11112), .Q(n6447) );
  CLKBU2 U197 ( .A(n6440), .Q(n11145) );
  NOR23 U198 ( .A(n11144), .B(n11099), .Q(n6449) );
  NOR23 U199 ( .A(n11144), .B(n11109), .Q(n6450) );
  NOR23 U200 ( .A(n11144), .B(n11107), .Q(n6451) );
  NOR23 U201 ( .A(n11144), .B(n11105), .Q(n6452) );
  NOR23 U202 ( .A(n11144), .B(n11102), .Q(n6453) );
  NOR23 U203 ( .A(n11144), .B(n11094), .Q(n6454) );
  NOR23 U204 ( .A(n11144), .B(n11141), .Q(n6455) );
  NOR23 U205 ( .A(n11144), .B(n11138), .Q(n6456) );
  CLKBU2 U206 ( .A(n6440), .Q(n11144) );
  NOR23 U207 ( .A(n11137), .B(n11133), .Q(n6457) );
  NOR23 U208 ( .A(n11137), .B(n11130), .Q(n6459) );
  NOR23 U209 ( .A(n11137), .B(n11127), .Q(n6461) );
  NOR23 U210 ( .A(n11137), .B(n11124), .Q(n6462) );
  NOR23 U211 ( .A(n11137), .B(n11121), .Q(n6463) );
  NOR23 U212 ( .A(n11137), .B(n11118), .Q(n6464) );
  NOR23 U213 ( .A(n11137), .B(n11115), .Q(n6465) );
  NOR23 U214 ( .A(n11137), .B(n11112), .Q(n6466) );
  CLKBU2 U215 ( .A(n6458), .Q(n11137) );
  NOR23 U216 ( .A(n11136), .B(n11099), .Q(n6467) );
  NOR23 U217 ( .A(n11136), .B(n11109), .Q(n6468) );
  NOR23 U218 ( .A(n11136), .B(n11107), .Q(n6469) );
  NOR23 U219 ( .A(n11136), .B(n11105), .Q(n6470) );
  NOR23 U220 ( .A(n11136), .B(n11102), .Q(n6472) );
  NOR23 U221 ( .A(n11136), .B(n11094), .Q(n6473) );
  NOR23 U222 ( .A(n11136), .B(n11141), .Q(n6474) );
  NOR23 U223 ( .A(n11136), .B(n11138), .Q(n6477) );
  CLKBU2 U224 ( .A(n6458), .Q(n11136) );
  NOR23 U225 ( .A(n11163), .B(n11135), .Q(n6275) );
  NOR23 U226 ( .A(n11163), .B(n11131), .Q(n6277) );
  NOR23 U227 ( .A(n11163), .B(n11128), .Q(n6279) );
  NOR23 U228 ( .A(n11163), .B(n11125), .Q(n6280) );
  NOR23 U229 ( .A(n11163), .B(n11122), .Q(n6281) );
  NOR23 U230 ( .A(n11163), .B(n11119), .Q(n6282) );
  NOR23 U231 ( .A(n11163), .B(n11116), .Q(n6283) );
  CLKBU2 U232 ( .A(n6215), .Q(n11116) );
  NOR23 U233 ( .A(n11163), .B(n11113), .Q(n6284) );
  CLKBU2 U234 ( .A(n6217), .Q(n11113) );
  NOR23 U235 ( .A(n11162), .B(n11101), .Q(n6285) );
  NOR23 U236 ( .A(n11162), .B(n11111), .Q(n6286) );
  NOR23 U237 ( .A(n11162), .B(n11108), .Q(n6287) );
  NOR23 U238 ( .A(n11162), .B(n11106), .Q(n6288) );
  NOR23 U239 ( .A(n11162), .B(n11103), .Q(n6290) );
  NOR23 U240 ( .A(n11162), .B(n11095), .Q(n6291) );
  NOR23 U241 ( .A(n11162), .B(n11143), .Q(n6292) );
  CLKBU2 U242 ( .A(n6196), .Q(n11143) );
  NOR23 U243 ( .A(n11162), .B(n11140), .Q(n6293) );
  CLKBU2 U244 ( .A(n6200), .Q(n11140) );
  NOR23 U245 ( .A(n11168), .B(n11134), .Q(n6201) );
  NOR23 U246 ( .A(n11168), .B(n11100), .Q(n6218) );
  NOR23 U247 ( .A(n11168), .B(n11110), .Q(n6220) );
  NOR23 U248 ( .A(n11168), .B(n11095), .Q(n6230) );
  NOR23 U249 ( .A(n11168), .B(n11142), .Q(n6232) );
  NOR23 U250 ( .A(n11168), .B(n11139), .Q(n6233) );
  CLKBU2 U251 ( .A(n6200), .Q(n11139) );
  NOR23 U252 ( .A(n11107), .B(n11092), .Q(n6494) );
  NOR23 U253 ( .A(n11105), .B(n11092), .Q(n6495) );
  NOR23 U254 ( .A(n11107), .B(n11169), .Q(n6224) );
  NOR23 U255 ( .A(n11105), .B(n11168), .Q(n6226) );
  CLKBU2 U256 ( .A(n6227), .Q(n11105) );
  NOR23 U257 ( .A(n11107), .B(n11098), .Q(n6223) );
  NOR23 U258 ( .A(n11105), .B(n11098), .Q(n6241) );
  NOR23 U259 ( .A(n11097), .B(n11099), .Q(n6194) );
  NOR23 U260 ( .A(n11097), .B(n11096), .Q(n6265) );
  NOR23 U261 ( .A(n11092), .B(n11094), .Q(n6193) );
  NOR23 U262 ( .A(n11102), .B(n11168), .Q(n6228) );
  NOR23 U263 ( .A(n11127), .B(n11097), .Q(n6418) );
  NOR23 U264 ( .A(n11124), .B(n11097), .Q(n6424) );
  NOR23 U265 ( .A(n11121), .B(n11097), .Q(n6435) );
  CLKBU2 U266 ( .A(n6211), .Q(n11121) );
  NOR23 U267 ( .A(n11118), .B(n11097), .Q(n6448) );
  CLKBU2 U268 ( .A(n6213), .Q(n11118) );
  NOR23 U269 ( .A(n11115), .B(n11097), .Q(n6460) );
  CLKBU2 U270 ( .A(n6215), .Q(n11115) );
  NOR23 U271 ( .A(n11112), .B(n11097), .Q(n6471) );
  CLKBU2 U272 ( .A(n6217), .Q(n11112) );
  NOR23 U273 ( .A(n11115), .B(n11092), .Q(n6489) );
  NOR23 U274 ( .A(n11112), .B(n11092), .Q(n6490) );
  NOR23 U275 ( .A(n11099), .B(n11092), .Q(n6491) );
  NOR23 U276 ( .A(n11109), .B(n11092), .Q(n6492) );
  CLKBU2 U277 ( .A(n6221), .Q(n11109) );
  NOR23 U278 ( .A(n11102), .B(n11092), .Q(n6496) );
  CLKBU2 U279 ( .A(n6229), .Q(n11102) );
  NOR23 U280 ( .A(n11130), .B(n11169), .Q(n6204) );
  NOR23 U281 ( .A(n11127), .B(n11169), .Q(n6206) );
  NOR23 U282 ( .A(n11124), .B(n11169), .Q(n6208) );
  NOR23 U283 ( .A(n11121), .B(n11169), .Q(n6210) );
  NOR23 U284 ( .A(n11118), .B(n11169), .Q(n6212) );
  NOR23 U285 ( .A(n11115), .B(n11169), .Q(n6214) );
  NOR23 U286 ( .A(n11112), .B(n11169), .Q(n6216) );
  NOR23 U287 ( .A(n11133), .B(n11093), .Q(n6479) );
  NOR23 U288 ( .A(n11130), .B(n11093), .Q(n6482) );
  NOR23 U289 ( .A(n11127), .B(n11093), .Q(n6484) );
  NOR23 U290 ( .A(n11124), .B(n11093), .Q(n6485) );
  NOR23 U291 ( .A(n11121), .B(n11093), .Q(n6486) );
  NOR23 U292 ( .A(n11118), .B(n11093), .Q(n6488) );
  NOR23 U293 ( .A(n11141), .B(n11093), .Q(n6195) );
  NOR23 U294 ( .A(n11138), .B(n11093), .Q(n6198) );
  NOR23 U295 ( .A(n11133), .B(n11098), .Q(n6416) );
  NOR23 U296 ( .A(n11130), .B(n11098), .Q(n6417) );
  NOR23 U297 ( .A(n11109), .B(n11098), .Q(n6199) );
  NOR23 U298 ( .A(n11102), .B(n11098), .Q(n6252) );
  NOR23 U299 ( .A(n11141), .B(n11098), .Q(n6278) );
  CLKBU2 U300 ( .A(n6196), .Q(n11141) );
  NOR23 U301 ( .A(n11138), .B(n11098), .Q(n6289) );
  CLKBU2 U302 ( .A(n6200), .Q(n11138) );
  BUF2 U303 ( .A(n6225), .Q(n11107) );
  BUF2 U304 ( .A(n6365), .Q(n11153) );
  BUF2 U305 ( .A(n6400), .Q(n11149) );
  BUF2 U306 ( .A(n6202), .Q(n11169) );
  BUF2 U307 ( .A(n6202), .Q(n11168) );
  BUF2 U308 ( .A(n6276), .Q(n11163) );
  BUF2 U309 ( .A(n6276), .Q(n11162) );
  BUF2 U310 ( .A(n6222), .Q(n11097) );
  BUF2 U315 ( .A(n6222), .Q(n11098) );
  BUF2 U320 ( .A(n6197), .Q(n11092) );
  BUF2 U325 ( .A(n6197), .Q(n11093) );
  INV3 U330 ( .A(n10863), .Q(n11315) );
  INV3 U331 ( .A(n10788), .Q(n11339) );
  INV3 U336 ( .A(n10871), .Q(n11318) );
  INV3 U341 ( .A(n10861), .Q(n11319) );
  INV3 U346 ( .A(n10856), .Q(n11316) );
  INV3 U351 ( .A(n10873), .Q(n11314) );
  INV3 U352 ( .A(n10876), .Q(n11317) );
  INV3 U357 ( .A(n10878), .Q(n11313) );
  INV3 U362 ( .A(n10851), .Q(n11320) );
  NOR21 U367 ( .A(n11321), .B(n11312), .Q(n10860) );
  NOR21 U372 ( .A(n11341), .B(n11332), .Q(n10709) );
  INV3 U373 ( .A(n10738), .Q(n11340) );
  INV3 U378 ( .A(n10732), .Q(n11326) );
  INV3 U383 ( .A(n10761), .Q(n11335) );
  INV3 U388 ( .A(n10810), .Q(n11334) );
  INV3 U393 ( .A(n10782), .Q(n11325) );
  INV3 U394 ( .A(n10708), .Q(n11331) );
  INV3 U395 ( .A(n10714), .Q(n11336) );
  INV3 U400 ( .A(n10685), .Q(n11327) );
  INV3 U405 ( .A(n10833), .Q(n11338) );
  INV3 U410 ( .A(n10827), .Q(n11324) );
  INV3 U415 ( .A(n10880), .Q(n11333) );
  INV3 U416 ( .A(n10842), .Q(n11337) );
  INV3 U421 ( .A(n10865), .Q(n11328) );
  INV3 U426 ( .A(n10805), .Q(n11329) );
  INV3 U431 ( .A(n10872), .Q(n11305) );
  INV3 U436 ( .A(n10862), .Q(n11306) );
  INV3 U437 ( .A(n10877), .Q(n11304) );
  INV3 U442 ( .A(n10879), .Q(n11308) );
  INV3 U447 ( .A(n10859), .Q(n11311) );
  INV3 U452 ( .A(n10854), .Q(n11307) );
  INV3 U457 ( .A(n10875), .Q(n11309) );
  NOR21 U458 ( .A(n11344), .B(waddr_1), .Q(n6483) );
  NOR21 U463 ( .A(waddr_1), .B(waddr_0), .Q(n6481) );
  NOR21 U468 ( .A(n11345), .B(waddr_0), .Q(n6475) );
  NOR21 U473 ( .A(n11347), .B(waddr_2), .Q(n6493) );
  NOR21 U478 ( .A(waddr_3), .B(waddr_2), .Q(n6480) );
  NOR21 U479 ( .A(n11346), .B(waddr_3), .Q(n6487) );
  NOR21 U480 ( .A(raddr_0), .B(raddr_1), .Q(n10858) );
  NOR21 U481 ( .A(raddr_4), .B(raddr_5), .Q(n10739) );
  NOR21 U486 ( .A(raddr_2), .B(raddr_3), .Q(n10864) );
  NOR21 U491 ( .A(raddr_6), .B(raddr_7), .Q(n10783) );
  BUF2 U496 ( .A(n6673), .Q(n10989) );
  BUF2 U501 ( .A(n6673), .Q(n10988) );
  BUF2 U502 ( .A(n11310), .Q(n6146) );
  BUF6 U507 ( .A(n6762), .Q(n11220) );
  BUF6 U512 ( .A(n6760), .Q(n11221) );
  BUF6 U517 ( .A(n6764), .Q(n11219) );
  BUF6 U522 ( .A(n6766), .Q(n11218) );
  BUF6 U523 ( .A(n6750), .Q(n11224) );
  BUF6 U528 ( .A(n6748), .Q(n11225) );
  BUF6 U533 ( .A(n6752), .Q(n11223) );
  BUF6 U538 ( .A(n6682), .Q(n11244) );
  BUF6 U543 ( .A(n6680), .Q(n11245) );
  BUF6 U544 ( .A(n6684), .Q(n11243) );
  BUF6 U549 ( .A(n6686), .Q(n11242) );
  BUF6 U554 ( .A(n6670), .Q(n11248) );
  BUF6 U559 ( .A(n6668), .Q(n11249) );
  BUF6 U564 ( .A(n6672), .Q(n11247) );
  BUF6 U565 ( .A(n6594), .Q(n11270) );
  BUF6 U566 ( .A(n6570), .Q(n11278) );
  BUF6 U571 ( .A(n6542), .Q(n11286) );
  BUF6 U576 ( .A(n6518), .Q(n11294) );
  BUF6 U581 ( .A(n6646), .Q(n11254) );
  BUF6 U586 ( .A(n6622), .Q(n11262) );
  BUF6 U587 ( .A(n6698), .Q(n11238) );
  BUF6 U592 ( .A(n6674), .Q(n11246) );
  BUF6 U597 ( .A(n6806), .Q(n11206) );
  BUF6 U602 ( .A(n6782), .Q(n11214) );
  BUF6 U607 ( .A(n6754), .Q(n11222) );
  BUF6 U608 ( .A(n6730), .Q(n11230) );
  BUF6 U613 ( .A(n6858), .Q(n11190) );
  BUF6 U618 ( .A(n6834), .Q(n11198) );
  BUF6 U623 ( .A(n6910), .Q(n11174) );
  BUF6 U628 ( .A(n6886), .Q(n11182) );
  BUF6 U629 ( .A(n6602), .Q(n11268) );
  BUF6 U634 ( .A(n6600), .Q(n11269) );
  BUF6 U639 ( .A(n6604), .Q(n11267) );
  BUF6 U644 ( .A(n6606), .Q(n11266) );
  BUF6 U649 ( .A(n6590), .Q(n11272) );
  BUF6 U650 ( .A(n6588), .Q(n11273) );
  BUF6 U651 ( .A(n6592), .Q(n11271) );
  BUF6 U652 ( .A(n6578), .Q(n11276) );
  BUF6 U657 ( .A(n6576), .Q(n11277) );
  BUF6 U662 ( .A(n6580), .Q(n11275) );
  BUF6 U667 ( .A(n6582), .Q(n11274) );
  BUF6 U672 ( .A(n6566), .Q(n11280) );
  BUF6 U673 ( .A(n6564), .Q(n11281) );
  BUF6 U678 ( .A(n6568), .Q(n11279) );
  BUF6 U683 ( .A(n6550), .Q(n11284) );
  BUF6 U688 ( .A(n6548), .Q(n11285) );
  BUF6 U693 ( .A(n6552), .Q(n11283) );
  BUF6 U694 ( .A(n6554), .Q(n11282) );
  BUF6 U699 ( .A(n6538), .Q(n11288) );
  BUF6 U704 ( .A(n6536), .Q(n11289) );
  BUF6 U709 ( .A(n6540), .Q(n11287) );
  BUF6 U714 ( .A(n6526), .Q(n11292) );
  BUF6 U715 ( .A(n6524), .Q(n11293) );
  BUF6 U720 ( .A(n6528), .Q(n11291) );
  BUF6 U725 ( .A(n6530), .Q(n11290) );
  BUF6 U730 ( .A(n6514), .Q(n11296) );
  BUF6 U735 ( .A(n6512), .Q(n11297) );
  BUF6 U736 ( .A(n6516), .Q(n11295) );
  BUF6 U737 ( .A(n6654), .Q(n11252) );
  BUF6 U742 ( .A(n6652), .Q(n11253) );
  BUF6 U747 ( .A(n6656), .Q(n11251) );
  BUF6 U752 ( .A(n6658), .Q(n11250) );
  BUF6 U757 ( .A(n6642), .Q(n11256) );
  BUF6 U758 ( .A(n6640), .Q(n11257) );
  BUF6 U763 ( .A(n6644), .Q(n11255) );
  BUF6 U768 ( .A(n6630), .Q(n11260) );
  BUF6 U773 ( .A(n6628), .Q(n11261) );
  BUF6 U778 ( .A(n6632), .Q(n11259) );
  BUF6 U779 ( .A(n6634), .Q(n11258) );
  BUF6 U784 ( .A(n6618), .Q(n11264) );
  BUF6 U789 ( .A(n6616), .Q(n11265) );
  BUF6 U794 ( .A(n6620), .Q(n11263) );
  BUF6 U799 ( .A(n6706), .Q(n11236) );
  BUF6 U800 ( .A(n6704), .Q(n11237) );
  BUF6 U805 ( .A(n6708), .Q(n11235) );
  BUF6 U810 ( .A(n6710), .Q(n11234) );
  BUF6 U815 ( .A(n6694), .Q(n11240) );
  BUF6 U820 ( .A(n6692), .Q(n11241) );
  BUF6 U821 ( .A(n6696), .Q(n11239) );
  BUF6 U822 ( .A(n6814), .Q(n11204) );
  BUF6 U823 ( .A(n6812), .Q(n11205) );
  BUF6 U828 ( .A(n6816), .Q(n11203) );
  BUF6 U833 ( .A(n6818), .Q(n11202) );
  BUF6 U838 ( .A(n6802), .Q(n11208) );
  BUF6 U843 ( .A(n6800), .Q(n11209) );
  BUF6 U844 ( .A(n6804), .Q(n11207) );
  BUF6 U849 ( .A(n6790), .Q(n11212) );
  BUF6 U854 ( .A(n6788), .Q(n11213) );
  BUF6 U859 ( .A(n6792), .Q(n11211) );
  BUF6 U864 ( .A(n6794), .Q(n11210) );
  BUF6 U865 ( .A(n6778), .Q(n11216) );
  BUF6 U870 ( .A(n6776), .Q(n11217) );
  BUF6 U875 ( .A(n6780), .Q(n11215) );
  BUF6 U880 ( .A(n6738), .Q(n11228) );
  BUF6 U885 ( .A(n6736), .Q(n11229) );
  BUF6 U886 ( .A(n6740), .Q(n11227) );
  BUF6 U891 ( .A(n6742), .Q(n11226) );
  BUF6 U896 ( .A(n6726), .Q(n11232) );
  BUF6 U901 ( .A(n6724), .Q(n11233) );
  BUF6 U906 ( .A(n6728), .Q(n11231) );
  BUF6 U907 ( .A(n6866), .Q(n11188) );
  BUF6 U908 ( .A(n6864), .Q(n11189) );
  BUF6 U913 ( .A(n6868), .Q(n11187) );
  BUF6 U918 ( .A(n6870), .Q(n11186) );
  BUF6 U923 ( .A(n6854), .Q(n11192) );
  BUF6 U928 ( .A(n6852), .Q(n11193) );
  BUF6 U929 ( .A(n6856), .Q(n11191) );
  BUF6 U934 ( .A(n6842), .Q(n11196) );
  BUF6 U939 ( .A(n6840), .Q(n11197) );
  BUF6 U944 ( .A(n6844), .Q(n11195) );
  BUF6 U949 ( .A(n6846), .Q(n11194) );
  BUF6 U950 ( .A(n6830), .Q(n11200) );
  BUF6 U955 ( .A(n6828), .Q(n11201) );
  BUF6 U960 ( .A(n6832), .Q(n11199) );
  BUF6 U965 ( .A(n6918), .Q(n11172) );
  BUF6 U970 ( .A(n6916), .Q(n11173) );
  BUF6 U971 ( .A(n6920), .Q(n11171) );
  BUF6 U976 ( .A(n6922), .Q(n11170) );
  BUF6 U981 ( .A(n6906), .Q(n11176) );
  BUF6 U986 ( .A(n6904), .Q(n11177) );
  BUF6 U991 ( .A(n6908), .Q(n11175) );
  BUF6 U992 ( .A(n6894), .Q(n11180) );
  BUF6 U993 ( .A(n6892), .Q(n11181) );
  BUF6 U994 ( .A(n6896), .Q(n11179) );
  BUF6 U999 ( .A(n6898), .Q(n11178) );
  BUF6 U1004 ( .A(n6882), .Q(n11184) );
  BUF6 U1009 ( .A(n6880), .Q(n11185) );
  BUF6 U1014 ( .A(n6884), .Q(n11183) );
  BUF2 U1015 ( .A(n11310), .Q(n6147) );
  BUF2 U1020 ( .A(n11310), .Q(n6145) );
  BUF2 U1025 ( .A(n6601), .Q(n11033) );
  BUF2 U1030 ( .A(n6599), .Q(n11035) );
  BUF2 U1035 ( .A(n6603), .Q(n11031) );
  BUF2 U1036 ( .A(n6605), .Q(n11029) );
  BUF2 U1041 ( .A(n6589), .Q(n11041) );
  BUF2 U1046 ( .A(n6587), .Q(n11043) );
  BUF2 U1051 ( .A(n6591), .Q(n11039) );
  BUF2 U1056 ( .A(n6577), .Q(n11049) );
  BUF2 U1057 ( .A(n6575), .Q(n11051) );
  BUF2 U1062 ( .A(n6579), .Q(n11047) );
  BUF2 U1067 ( .A(n6581), .Q(n11045) );
  BUF2 U1072 ( .A(n6565), .Q(n11057) );
  BUF2 U1077 ( .A(n6563), .Q(n11059) );
  BUF2 U1078 ( .A(n6567), .Q(n11055) );
  BUF2 U1079 ( .A(n6549), .Q(n11065) );
  BUF2 U1084 ( .A(n6547), .Q(n11067) );
  BUF2 U1089 ( .A(n6551), .Q(n11063) );
  BUF2 U1094 ( .A(n6553), .Q(n11061) );
  BUF2 U1099 ( .A(n6537), .Q(n11073) );
  BUF2 U1100 ( .A(n6535), .Q(n11075) );
  BUF2 U1105 ( .A(n6539), .Q(n11071) );
  BUF2 U1110 ( .A(n6525), .Q(n11081) );
  BUF2 U1115 ( .A(n6523), .Q(n11083) );
  BUF2 U1120 ( .A(n6527), .Q(n11079) );
  BUF2 U1121 ( .A(n6529), .Q(n11077) );
  BUF2 U1126 ( .A(n6513), .Q(n11089) );
  BUF2 U1131 ( .A(n6511), .Q(n11091) );
  BUF2 U1136 ( .A(n6515), .Q(n11087) );
  BUF2 U1141 ( .A(n6653), .Q(n11001) );
  BUF2 U1142 ( .A(n6651), .Q(n11003) );
  BUF2 U1147 ( .A(n6655), .Q(n10999) );
  BUF2 U1152 ( .A(n6657), .Q(n10997) );
  BUF2 U1157 ( .A(n6641), .Q(n11009) );
  BUF2 U1162 ( .A(n6639), .Q(n11011) );
  BUF2 U1163 ( .A(n6643), .Q(n11007) );
  BUF2 U1164 ( .A(n6629), .Q(n11017) );
  BUF2 U1165 ( .A(n6627), .Q(n11019) );
  BUF2 U1170 ( .A(n6631), .Q(n11015) );
  BUF2 U1175 ( .A(n6633), .Q(n11013) );
  BUF2 U1180 ( .A(n6617), .Q(n11025) );
  BUF2 U1185 ( .A(n6615), .Q(n11027) );
  BUF2 U1186 ( .A(n6619), .Q(n11023) );
  BUF2 U1191 ( .A(n6705), .Q(n10969) );
  BUF2 U1196 ( .A(n6703), .Q(n10971) );
  BUF2 U1201 ( .A(n6707), .Q(n10967) );
  BUF2 U1206 ( .A(n6709), .Q(n10965) );
  BUF2 U1207 ( .A(n6693), .Q(n10977) );
  BUF2 U1212 ( .A(n6691), .Q(n10979) );
  BUF2 U1217 ( .A(n6695), .Q(n10975) );
  BUF2 U1222 ( .A(n6813), .Q(n10905) );
  BUF2 U1227 ( .A(n6811), .Q(n10907) );
  BUF2 U1228 ( .A(n6815), .Q(n10903) );
  BUF2 U1233 ( .A(n6817), .Q(n10901) );
  BUF2 U1238 ( .A(n6801), .Q(n10913) );
  BUF2 U1243 ( .A(n6799), .Q(n10915) );
  BUF2 U1248 ( .A(n6803), .Q(n10911) );
  BUF2 U1249 ( .A(n6789), .Q(n10921) );
  BUF2 U1250 ( .A(n6787), .Q(n10923) );
  BUF2 U1255 ( .A(n6791), .Q(n10919) );
  BUF2 U1260 ( .A(n6793), .Q(n10917) );
  BUF2 U1265 ( .A(n6777), .Q(n10929) );
  BUF2 U1270 ( .A(n6775), .Q(n10931) );
  BUF2 U1271 ( .A(n6779), .Q(n10927) );
  BUF2 U1276 ( .A(n6737), .Q(n10953) );
  BUF2 U1281 ( .A(n6735), .Q(n10955) );
  BUF2 U1286 ( .A(n6739), .Q(n10951) );
  BUF2 U1291 ( .A(n6741), .Q(n10949) );
  BUF2 U1292 ( .A(n6725), .Q(n10961) );
  BUF2 U1297 ( .A(n6723), .Q(n10963) );
  BUF2 U1302 ( .A(n6727), .Q(n10959) );
  BUF2 U1307 ( .A(n6865), .Q(n6185) );
  BUF2 U1312 ( .A(n6863), .Q(n6187) );
  BUF2 U1313 ( .A(n6867), .Q(n6183) );
  BUF2 U1318 ( .A(n6869), .Q(n6181) );
  BUF2 U1323 ( .A(n6853), .Q(n10881) );
  BUF2 U1328 ( .A(n6851), .Q(n10883) );
  BUF2 U1333 ( .A(n6855), .Q(n6191) );
  BUF2 U1334 ( .A(n6841), .Q(n10889) );
  BUF2 U1335 ( .A(n6839), .Q(n10891) );
  BUF2 U1336 ( .A(n6843), .Q(n10887) );
  BUF2 U1341 ( .A(n6845), .Q(n10885) );
  BUF2 U1346 ( .A(n6829), .Q(n10897) );
  BUF2 U1351 ( .A(n6827), .Q(n10899) );
  BUF2 U1356 ( .A(n6831), .Q(n10895) );
  BUF2 U1357 ( .A(n6917), .Q(n6153) );
  BUF2 U1362 ( .A(n6915), .Q(n6155) );
  BUF2 U1367 ( .A(n6919), .Q(n6151) );
  BUF2 U1372 ( .A(n6921), .Q(n6149) );
  BUF2 U1377 ( .A(n6905), .Q(n6161) );
  BUF2 U1378 ( .A(n6903), .Q(n6163) );
  BUF2 U1383 ( .A(n6907), .Q(n6159) );
  BUF2 U1388 ( .A(n6893), .Q(n6169) );
  BUF2 U1393 ( .A(n6891), .Q(n6171) );
  BUF2 U1398 ( .A(n6895), .Q(n6167) );
  BUF2 U1399 ( .A(n6897), .Q(n6165) );
  BUF2 U1404 ( .A(n6881), .Q(n6177) );
  BUF2 U1409 ( .A(n6879), .Q(n6179) );
  BUF2 U1414 ( .A(n6883), .Q(n6175) );
  BUF2 U1419 ( .A(n6601), .Q(n11032) );
  BUF2 U1420 ( .A(n6599), .Q(n11034) );
  BUF2 U1421 ( .A(n6603), .Q(n11030) );
  BUF2 U1426 ( .A(n6605), .Q(n11028) );
  BUF2 U1431 ( .A(n6589), .Q(n11040) );
  BUF2 U1436 ( .A(n6587), .Q(n11042) );
  BUF2 U1441 ( .A(n6591), .Q(n11038) );
  BUF2 U1442 ( .A(n6577), .Q(n11048) );
  BUF2 U1447 ( .A(n6575), .Q(n11050) );
  BUF2 U1452 ( .A(n6579), .Q(n11046) );
  BUF2 U1457 ( .A(n6581), .Q(n11044) );
  BUF2 U1462 ( .A(n6565), .Q(n11056) );
  BUF2 U1463 ( .A(n6563), .Q(n11058) );
  BUF2 U1468 ( .A(n6567), .Q(n11054) );
  BUF2 U1473 ( .A(n6549), .Q(n11064) );
  BUF2 U1478 ( .A(n6547), .Q(n11066) );
  BUF2 U1483 ( .A(n6551), .Q(n11062) );
  BUF2 U1484 ( .A(n6553), .Q(n11060) );
  BUF2 U1489 ( .A(n6537), .Q(n11072) );
  BUF2 U1494 ( .A(n6535), .Q(n11074) );
  BUF2 U1499 ( .A(n6539), .Q(n11070) );
  BUF2 U1504 ( .A(n6525), .Q(n11080) );
  BUF2 U1505 ( .A(n6523), .Q(n11082) );
  BUF2 U1506 ( .A(n6527), .Q(n11078) );
  BUF2 U1507 ( .A(n6529), .Q(n11076) );
  BUF2 U1512 ( .A(n6513), .Q(n11088) );
  BUF2 U1517 ( .A(n6511), .Q(n11090) );
  BUF2 U1522 ( .A(n6515), .Q(n11086) );
  BUF2 U1527 ( .A(n6653), .Q(n11000) );
  BUF2 U1528 ( .A(n6651), .Q(n11002) );
  BUF2 U1533 ( .A(n6655), .Q(n10998) );
  BUF2 U1538 ( .A(n6657), .Q(n10996) );
  BUF2 U1543 ( .A(n6641), .Q(n11008) );
  BUF2 U1548 ( .A(n6639), .Q(n11010) );
  BUF2 U1549 ( .A(n6643), .Q(n11006) );
  BUF2 U1554 ( .A(n6629), .Q(n11016) );
  BUF2 U1559 ( .A(n6627), .Q(n11018) );
  BUF2 U1564 ( .A(n6631), .Q(n11014) );
  BUF2 U1569 ( .A(n6633), .Q(n11012) );
  BUF2 U1570 ( .A(n6617), .Q(n11024) );
  BUF2 U1575 ( .A(n6615), .Q(n11026) );
  BUF2 U1580 ( .A(n6619), .Q(n11022) );
  BUF2 U1585 ( .A(n6705), .Q(n10968) );
  BUF2 U1590 ( .A(n6703), .Q(n10970) );
  BUF2 U1591 ( .A(n6707), .Q(n10966) );
  BUF2 U1592 ( .A(n6709), .Q(n10964) );
  BUF2 U1597 ( .A(n6693), .Q(n10976) );
  BUF2 U1602 ( .A(n6691), .Q(n10978) );
  BUF2 U1607 ( .A(n6695), .Q(n10974) );
  BUF2 U1612 ( .A(n6813), .Q(n10904) );
  BUF2 U1613 ( .A(n6811), .Q(n10906) );
  BUF2 U1618 ( .A(n6815), .Q(n10902) );
  BUF2 U1623 ( .A(n6817), .Q(n10900) );
  BUF2 U1628 ( .A(n6801), .Q(n10912) );
  BUF2 U1633 ( .A(n6799), .Q(n10914) );
  BUF2 U1634 ( .A(n6803), .Q(n10910) );
  BUF2 U1639 ( .A(n6789), .Q(n10920) );
  BUF2 U1644 ( .A(n6787), .Q(n10922) );
  BUF2 U1649 ( .A(n6791), .Q(n10918) );
  BUF2 U1654 ( .A(n6793), .Q(n10916) );
  BUF2 U1655 ( .A(n6777), .Q(n10928) );
  BUF2 U1660 ( .A(n6775), .Q(n10930) );
  BUF2 U1665 ( .A(n6779), .Q(n10926) );
  BUF2 U1670 ( .A(n6737), .Q(n10952) );
  BUF2 U1675 ( .A(n6735), .Q(n10954) );
  BUF2 U1676 ( .A(n6739), .Q(n10950) );
  BUF2 U1677 ( .A(n6741), .Q(n10948) );
  BUF2 U1678 ( .A(n6725), .Q(n10960) );
  BUF2 U1683 ( .A(n6723), .Q(n10962) );
  BUF2 U1688 ( .A(n6727), .Q(n10958) );
  BUF2 U1693 ( .A(n6865), .Q(n6184) );
  BUF2 U1698 ( .A(n6863), .Q(n6186) );
  BUF2 U1699 ( .A(n6867), .Q(n6182) );
  BUF2 U1704 ( .A(n6869), .Q(n6180) );
  BUF2 U1709 ( .A(n6853), .Q(n6192) );
  BUF2 U1714 ( .A(n6851), .Q(n10882) );
  BUF2 U1719 ( .A(n6855), .Q(n6190) );
  BUF2 U1720 ( .A(n6841), .Q(n10888) );
  BUF2 U1725 ( .A(n6839), .Q(n10890) );
  BUF2 U1730 ( .A(n6843), .Q(n10886) );
  BUF2 U1735 ( .A(n6845), .Q(n10884) );
  BUF2 U1740 ( .A(n6829), .Q(n10896) );
  BUF2 U1741 ( .A(n6827), .Q(n10898) );
  BUF2 U1746 ( .A(n6831), .Q(n10894) );
  BUF2 U1751 ( .A(n6917), .Q(n6152) );
  BUF2 U1756 ( .A(n6915), .Q(n6154) );
  BUF2 U1761 ( .A(n6919), .Q(n6150) );
  BUF2 U1762 ( .A(n6921), .Q(n6148) );
  BUF2 U1763 ( .A(n6905), .Q(n6160) );
  BUF2 U1768 ( .A(n6903), .Q(n6162) );
  BUF2 U1773 ( .A(n6907), .Q(n6158) );
  BUF2 U1778 ( .A(n6893), .Q(n6168) );
  BUF2 U1783 ( .A(n6891), .Q(n6170) );
  BUF2 U1784 ( .A(n6895), .Q(n6166) );
  BUF2 U1789 ( .A(n6897), .Q(n6164) );
  BUF2 U1794 ( .A(n6881), .Q(n6176) );
  BUF2 U1799 ( .A(n6879), .Q(n6178) );
  BUF2 U1804 ( .A(n6883), .Q(n6174) );
  BUF2 U1805 ( .A(n6761), .Q(n10937) );
  BUF2 U1810 ( .A(n6759), .Q(n10939) );
  BUF2 U1815 ( .A(n6763), .Q(n10935) );
  BUF2 U1820 ( .A(n6765), .Q(n10933) );
  BUF2 U1825 ( .A(n6749), .Q(n10945) );
  BUF2 U1826 ( .A(n6747), .Q(n10947) );
  BUF2 U1831 ( .A(n6751), .Q(n10943) );
  BUF2 U1836 ( .A(n6753), .Q(n10941) );
  BUF2 U1841 ( .A(n6761), .Q(n10936) );
  BUF2 U1846 ( .A(n6759), .Q(n10938) );
  BUF2 U1847 ( .A(n6763), .Q(n10934) );
  BUF2 U1848 ( .A(n6765), .Q(n10932) );
  BUF2 U1849 ( .A(n6749), .Q(n10944) );
  BUF2 U1854 ( .A(n6747), .Q(n10946) );
  BUF2 U1859 ( .A(n6751), .Q(n10942) );
  BUF2 U1864 ( .A(n6753), .Q(n10940) );
  BUF2 U1869 ( .A(n6681), .Q(n10985) );
  BUF2 U1870 ( .A(n6679), .Q(n10987) );
  BUF2 U1875 ( .A(n6683), .Q(n10983) );
  BUF2 U1880 ( .A(n6685), .Q(n10981) );
  BUF2 U1885 ( .A(n6669), .Q(n10993) );
  BUF2 U1890 ( .A(n6667), .Q(n10995) );
  BUF2 U1891 ( .A(n6671), .Q(n10991) );
  BUF2 U1896 ( .A(n6681), .Q(n10984) );
  BUF2 U1901 ( .A(n6679), .Q(n10986) );
  BUF2 U1906 ( .A(n6683), .Q(n10982) );
  BUF2 U1911 ( .A(n6685), .Q(n10980) );
  BUF2 U1912 ( .A(n6669), .Q(n10992) );
  BUF2 U1917 ( .A(n6667), .Q(n10994) );
  BUF2 U1922 ( .A(n6671), .Q(n10990) );
  BUF2 U1927 ( .A(n6593), .Q(n11037) );
  BUF2 U1932 ( .A(n6541), .Q(n11069) );
  BUF2 U1933 ( .A(n6645), .Q(n11005) );
  BUF2 U1934 ( .A(n6697), .Q(n10973) );
  BUF2 U1939 ( .A(n6781), .Q(n10925) );
  BUF2 U1944 ( .A(n6593), .Q(n11036) );
  BUF2 U1949 ( .A(n6541), .Q(n11068) );
  BUF2 U1954 ( .A(n6645), .Q(n11004) );
  BUF2 U1955 ( .A(n6697), .Q(n10972) );
  BUF2 U1960 ( .A(n6781), .Q(n10924) );
  BUF2 U1965 ( .A(n6569), .Q(n11053) );
  BUF2 U1970 ( .A(n6517), .Q(n11085) );
  BUF2 U1975 ( .A(n6621), .Q(n11021) );
  BUF2 U1976 ( .A(n6805), .Q(n10909) );
  BUF2 U1981 ( .A(n6729), .Q(n10957) );
  BUF2 U1986 ( .A(n6857), .Q(n6189) );
  BUF2 U1991 ( .A(n6833), .Q(n10893) );
  BUF2 U1996 ( .A(n6909), .Q(n6157) );
  BUF2 U1997 ( .A(n6885), .Q(n6173) );
  BUF2 U2002 ( .A(n6569), .Q(n11052) );
  BUF2 U2007 ( .A(n6517), .Q(n11084) );
  BUF2 U2012 ( .A(n6621), .Q(n11020) );
  BUF2 U2017 ( .A(n6805), .Q(n10908) );
  BUF2 U2018 ( .A(n6729), .Q(n10956) );
  BUF2 U2019 ( .A(n6857), .Q(n6188) );
  BUF2 U2020 ( .A(n6833), .Q(n10892) );
  BUF2 U2025 ( .A(n6909), .Q(n6156) );
  BUF2 U2030 ( .A(n6885), .Q(n6172) );
  NAND22 U2035 ( .A(n11330), .B(n6147), .Q(n6673) );
  NAND22 U2040 ( .A(n6478), .B(n6476), .Q(n6200) );
  BUF2 U2041 ( .A(n6211), .Q(n11122) );
  BUF2 U2046 ( .A(n6203), .Q(n11134) );
  BUF2 U2051 ( .A(n6219), .Q(n11100) );
  BUF2 U2056 ( .A(n6205), .Q(n11131) );
  BUF2 U2061 ( .A(n6221), .Q(n11110) );
  BUF2 U2062 ( .A(n6207), .Q(n11128) );
  BUF2 U2067 ( .A(n6229), .Q(n11103) );
  BUF2 U2072 ( .A(n6209), .Q(n11125) );
  BUF2 U2077 ( .A(n6205), .Q(n11130) );
  BUF2 U2082 ( .A(n6207), .Q(n11127) );
  BUF2 U2083 ( .A(n6209), .Q(n11124) );
  BUF2 U2088 ( .A(n6203), .Q(n11133) );
  BUF2 U2093 ( .A(n6219), .Q(n11099) );
  BUF2 U2098 ( .A(n6203), .Q(n11135) );
  BUF2 U2103 ( .A(n6219), .Q(n11101) );
  BUF2 U2104 ( .A(n6211), .Q(n11123) );
  BUF2 U2105 ( .A(n6231), .Q(n11095) );
  BUF2 U2110 ( .A(n6221), .Q(n11111) );
  BUF2 U2115 ( .A(n6205), .Q(n11132) );
  BUF2 U2120 ( .A(n6213), .Q(n11120) );
  BUF2 U2125 ( .A(n6231), .Q(n11096) );
  BUF2 U2126 ( .A(n6207), .Q(n11129) );
  BUF2 U2131 ( .A(n6229), .Q(n11104) );
  BUF2 U2136 ( .A(n6209), .Q(n11126) );
  INV3 U2141 ( .A(n10756), .Q(n11330) );
  NAND22 U2146 ( .A(n10733), .B(n10709), .Q(n10756) );
  NAND22 U2147 ( .A(n11314), .B(n11339), .Q(n6762) );
  NAND22 U2152 ( .A(n11318), .B(n11339), .Q(n6760) );
  NAND22 U2157 ( .A(n11317), .B(n11339), .Q(n6764) );
  NAND22 U2162 ( .A(n11313), .B(n11339), .Q(n6766) );
  NAND22 U2167 ( .A(n11316), .B(n11339), .Q(n6750) );
  NAND22 U2168 ( .A(n11320), .B(n11339), .Q(n6748) );
  NAND22 U2173 ( .A(n11319), .B(n11339), .Q(n6752) );
  NAND22 U2178 ( .A(n11314), .B(n11330), .Q(n6682) );
  NAND22 U2183 ( .A(n11318), .B(n11330), .Q(n6680) );
  NAND22 U2188 ( .A(n11317), .B(n11330), .Q(n6684) );
  NAND22 U2189 ( .A(n11313), .B(n11330), .Q(n6686) );
  NAND22 U2190 ( .A(n11316), .B(n11330), .Q(n6670) );
  NAND22 U2191 ( .A(n11320), .B(n11330), .Q(n6668) );
  NAND22 U2196 ( .A(n11319), .B(n11330), .Q(n6672) );
  NAND22 U2201 ( .A(n11331), .B(n11315), .Q(n6594) );
  NAND22 U2206 ( .A(n11340), .B(n11315), .Q(n6570) );
  NAND22 U2211 ( .A(n11327), .B(n11315), .Q(n6542) );
  NAND22 U2212 ( .A(n11336), .B(n11315), .Q(n6518) );
  NAND22 U2217 ( .A(n11326), .B(n11315), .Q(n6646) );
  NAND22 U2222 ( .A(n11335), .B(n11315), .Q(n6622) );
  NAND22 U2227 ( .A(n11330), .B(n11315), .Q(n6698) );
  NAND22 U2232 ( .A(n11339), .B(n11315), .Q(n6674) );
  NAND22 U2233 ( .A(n11329), .B(n11315), .Q(n6806) );
  NAND22 U2238 ( .A(n11338), .B(n11315), .Q(n6782) );
  NAND22 U2243 ( .A(n11325), .B(n11315), .Q(n6754) );
  NAND22 U2248 ( .A(n11334), .B(n11315), .Q(n6730) );
  NAND22 U2253 ( .A(n11324), .B(n11315), .Q(n6858) );
  NAND22 U2254 ( .A(n11333), .B(n11315), .Q(n6834) );
  NAND22 U2259 ( .A(n11328), .B(n11315), .Q(n6910) );
  NAND22 U2264 ( .A(n11337), .B(n11315), .Q(n6886) );
  NAND22 U2269 ( .A(n11336), .B(n11314), .Q(n6602) );
  NAND22 U2274 ( .A(n11336), .B(n11313), .Q(n6606) );
  NAND22 U2275 ( .A(n11336), .B(n11316), .Q(n6590) );
  NAND22 U2276 ( .A(n11331), .B(n11314), .Q(n6578) );
  NAND22 U2281 ( .A(n11331), .B(n11313), .Q(n6582) );
  NAND22 U2286 ( .A(n11331), .B(n11316), .Q(n6566) );
  NAND22 U2291 ( .A(n11337), .B(n11314), .Q(n6550) );
  NAND22 U2296 ( .A(n11337), .B(n11313), .Q(n6554) );
  NAND22 U2297 ( .A(n11337), .B(n11316), .Q(n6538) );
  NAND22 U2302 ( .A(n11327), .B(n11314), .Q(n6526) );
  NAND22 U2307 ( .A(n11327), .B(n11313), .Q(n6530) );
  NAND22 U2312 ( .A(n11327), .B(n11316), .Q(n6514) );
  NAND22 U2317 ( .A(n11340), .B(n11314), .Q(n6654) );
  NAND22 U2318 ( .A(n11340), .B(n11313), .Q(n6658) );
  NAND22 U2323 ( .A(n11340), .B(n11316), .Q(n6642) );
  NAND22 U2328 ( .A(n11326), .B(n11314), .Q(n6630) );
  NAND22 U2333 ( .A(n11326), .B(n11313), .Q(n6634) );
  NAND22 U2338 ( .A(n11326), .B(n11316), .Q(n6618) );
  NAND22 U2339 ( .A(n11335), .B(n11314), .Q(n6706) );
  NAND22 U2344 ( .A(n11335), .B(n11313), .Q(n6710) );
  NAND22 U2349 ( .A(n11335), .B(n11316), .Q(n6694) );
  NAND22 U2354 ( .A(n11334), .B(n11314), .Q(n6814) );
  NAND22 U2359 ( .A(n11334), .B(n11313), .Q(n6818) );
  NAND22 U2360 ( .A(n11334), .B(n11316), .Q(n6802) );
  NAND22 U2361 ( .A(n11329), .B(n11314), .Q(n6790) );
  NAND22 U2362 ( .A(n11329), .B(n11313), .Q(n6794) );
  NAND22 U2367 ( .A(n11329), .B(n11316), .Q(n6778) );
  NAND22 U2372 ( .A(n11325), .B(n11314), .Q(n6738) );
  NAND22 U2377 ( .A(n11325), .B(n11313), .Q(n6742) );
  NAND22 U2382 ( .A(n11325), .B(n11316), .Q(n6726) );
  NAND22 U2383 ( .A(n11338), .B(n11314), .Q(n6866) );
  NAND22 U2388 ( .A(n11338), .B(n11313), .Q(n6870) );
  NAND22 U2393 ( .A(n11338), .B(n11316), .Q(n6854) );
  NAND22 U2398 ( .A(n11324), .B(n11314), .Q(n6842) );
  NAND22 U2403 ( .A(n11324), .B(n11313), .Q(n6846) );
  NAND22 U2404 ( .A(n11324), .B(n11316), .Q(n6830) );
  NAND22 U2409 ( .A(n11333), .B(n11314), .Q(n6918) );
  NAND22 U2414 ( .A(n11333), .B(n11313), .Q(n6922) );
  NAND22 U2419 ( .A(n11333), .B(n11316), .Q(n6906) );
  NAND22 U2424 ( .A(n11328), .B(n11314), .Q(n6894) );
  NAND22 U2425 ( .A(n11328), .B(n11313), .Q(n6898) );
  NAND22 U2430 ( .A(n11328), .B(n11316), .Q(n6882) );
  NAND22 U2435 ( .A(n11336), .B(n11318), .Q(n6600) );
  NAND22 U2440 ( .A(n11331), .B(n11318), .Q(n6576) );
  NAND22 U2445 ( .A(n11337), .B(n11318), .Q(n6548) );
  NAND22 U2446 ( .A(n11327), .B(n11318), .Q(n6524) );
  NAND22 U2447 ( .A(n11340), .B(n11318), .Q(n6652) );
  NAND22 U2452 ( .A(n11326), .B(n11318), .Q(n6628) );
  NAND22 U2457 ( .A(n11335), .B(n11318), .Q(n6704) );
  NAND22 U2462 ( .A(n11334), .B(n11318), .Q(n6812) );
  NAND22 U2467 ( .A(n11329), .B(n11318), .Q(n6788) );
  NAND22 U2468 ( .A(n11325), .B(n11318), .Q(n6736) );
  NAND22 U2473 ( .A(n11338), .B(n11318), .Q(n6864) );
  NAND22 U2478 ( .A(n11324), .B(n11318), .Q(n6840) );
  NAND22 U2483 ( .A(n11333), .B(n11318), .Q(n6916) );
  NAND22 U2488 ( .A(n11328), .B(n11318), .Q(n6892) );
  NAND22 U2489 ( .A(n11336), .B(n11317), .Q(n6604) );
  NAND22 U2494 ( .A(n11336), .B(n11320), .Q(n6588) );
  NAND22 U2499 ( .A(n11331), .B(n11317), .Q(n6580) );
  NAND22 U2504 ( .A(n11331), .B(n11320), .Q(n6564) );
  NAND22 U2509 ( .A(n11337), .B(n11317), .Q(n6552) );
  NAND22 U2510 ( .A(n11337), .B(n11320), .Q(n6536) );
  NAND22 U2515 ( .A(n11327), .B(n11317), .Q(n6528) );
  NAND22 U2520 ( .A(n11327), .B(n11320), .Q(n6512) );
  NAND22 U2525 ( .A(n11340), .B(n11317), .Q(n6656) );
  NAND22 U2530 ( .A(n11340), .B(n11320), .Q(n6640) );
  NAND22 U2531 ( .A(n11326), .B(n11317), .Q(n6632) );
  NAND22 U2532 ( .A(n11326), .B(n11320), .Q(n6616) );
  NAND22 U2533 ( .A(n11335), .B(n11317), .Q(n6708) );
  NAND22 U2538 ( .A(n11335), .B(n11320), .Q(n6692) );
  NAND22 U2543 ( .A(n11334), .B(n11317), .Q(n6816) );
  NAND22 U2548 ( .A(n11334), .B(n11320), .Q(n6800) );
  NAND22 U2553 ( .A(n11329), .B(n11317), .Q(n6792) );
  NAND22 U2554 ( .A(n11329), .B(n11320), .Q(n6776) );
  NAND22 U2559 ( .A(n11325), .B(n11317), .Q(n6740) );
  NAND22 U2564 ( .A(n11325), .B(n11320), .Q(n6724) );
  NAND22 U2569 ( .A(n11338), .B(n11317), .Q(n6868) );
  NAND22 U2574 ( .A(n11338), .B(n11320), .Q(n6852) );
  NAND22 U2575 ( .A(n11324), .B(n11317), .Q(n6844) );
  NAND22 U2580 ( .A(n11324), .B(n11320), .Q(n6828) );
  NAND22 U2585 ( .A(n11333), .B(n11317), .Q(n6920) );
  NAND22 U2590 ( .A(n11333), .B(n11320), .Q(n6904) );
  NAND22 U2595 ( .A(n11328), .B(n11317), .Q(n6896) );
  NAND22 U2596 ( .A(n11328), .B(n11320), .Q(n6880) );
  NAND22 U2601 ( .A(n11336), .B(n11319), .Q(n6592) );
  NAND22 U2606 ( .A(n11331), .B(n11319), .Q(n6568) );
  NAND22 U2611 ( .A(n11337), .B(n11319), .Q(n6540) );
  NAND22 U2616 ( .A(n11327), .B(n11319), .Q(n6516) );
  NAND22 U2617 ( .A(n11340), .B(n11319), .Q(n6644) );
  NAND22 U2618 ( .A(n11326), .B(n11319), .Q(n6620) );
  NAND22 U2623 ( .A(n11335), .B(n11319), .Q(n6696) );
  NAND22 U2628 ( .A(n11334), .B(n11319), .Q(n6804) );
  NAND22 U2633 ( .A(n11329), .B(n11319), .Q(n6780) );
  NAND22 U2638 ( .A(n11325), .B(n11319), .Q(n6728) );
  NAND22 U2639 ( .A(n11338), .B(n11319), .Q(n6856) );
  NAND22 U2644 ( .A(n11324), .B(n11319), .Q(n6832) );
  NAND22 U2649 ( .A(n11333), .B(n11319), .Q(n6908) );
  NAND22 U2654 ( .A(n11328), .B(n11319), .Q(n6884) );
  NAND22 U2659 ( .A(n11336), .B(n11309), .Q(n6601) );
  NAND22 U2660 ( .A(n11336), .B(n11305), .Q(n6599) );
  NAND22 U2665 ( .A(n11331), .B(n11309), .Q(n6577) );
  NAND22 U2670 ( .A(n11331), .B(n11305), .Q(n6575) );
  NAND22 U2675 ( .A(n11337), .B(n11309), .Q(n6549) );
  NAND22 U2680 ( .A(n11337), .B(n11305), .Q(n6547) );
  NAND22 U2681 ( .A(n11327), .B(n11309), .Q(n6525) );
  NAND22 U2686 ( .A(n11327), .B(n11305), .Q(n6523) );
  NAND22 U2691 ( .A(n11340), .B(n11309), .Q(n6653) );
  NAND22 U2696 ( .A(n11340), .B(n11305), .Q(n6651) );
  NAND22 U2701 ( .A(n11326), .B(n11309), .Q(n6629) );
  NAND22 U2702 ( .A(n11326), .B(n11305), .Q(n6627) );
  NAND22 U2703 ( .A(n11335), .B(n11309), .Q(n6705) );
  NAND22 U2704 ( .A(n11335), .B(n11305), .Q(n6703) );
  NAND22 U2709 ( .A(n11334), .B(n11309), .Q(n6813) );
  NAND22 U2714 ( .A(n11334), .B(n11305), .Q(n6811) );
  NAND22 U2719 ( .A(n11329), .B(n11309), .Q(n6789) );
  NAND22 U2724 ( .A(n11329), .B(n11305), .Q(n6787) );
  NAND22 U2725 ( .A(n11325), .B(n11309), .Q(n6737) );
  NAND22 U2730 ( .A(n11325), .B(n11305), .Q(n6735) );
  NAND22 U2735 ( .A(n11338), .B(n11309), .Q(n6865) );
  NAND22 U2740 ( .A(n11338), .B(n11305), .Q(n6863) );
  NAND22 U2745 ( .A(n11324), .B(n11309), .Q(n6841) );
  NAND22 U2746 ( .A(n11324), .B(n11305), .Q(n6839) );
  NAND22 U2751 ( .A(n11333), .B(n11309), .Q(n6917) );
  NAND22 U2756 ( .A(n11333), .B(n11305), .Q(n6915) );
  NAND22 U2761 ( .A(n11328), .B(n11309), .Q(n6893) );
  NAND22 U2766 ( .A(n11328), .B(n11305), .Q(n6891) );
  NAND22 U2767 ( .A(n11336), .B(n11304), .Q(n6603) );
  NAND22 U2772 ( .A(n11336), .B(n11307), .Q(n6587) );
  NAND22 U2777 ( .A(n11331), .B(n11304), .Q(n6579) );
  NAND22 U2782 ( .A(n11331), .B(n11307), .Q(n6563) );
  NAND22 U2787 ( .A(n11337), .B(n11304), .Q(n6551) );
  NAND22 U2788 ( .A(n11337), .B(n11307), .Q(n6535) );
  NAND22 U2789 ( .A(n11327), .B(n11304), .Q(n6527) );
  NAND22 U2794 ( .A(n11327), .B(n11307), .Q(n6511) );
  NAND22 U2799 ( .A(n11340), .B(n11304), .Q(n6655) );
  NAND22 U2804 ( .A(n11340), .B(n11307), .Q(n6639) );
  NAND22 U2809 ( .A(n11326), .B(n11304), .Q(n6631) );
  NAND22 U2810 ( .A(n11326), .B(n11307), .Q(n6615) );
  NAND22 U2815 ( .A(n11335), .B(n11304), .Q(n6707) );
  NAND22 U2820 ( .A(n11335), .B(n11307), .Q(n6691) );
  NAND22 U2825 ( .A(n11334), .B(n11304), .Q(n6815) );
  NAND22 U2830 ( .A(n11334), .B(n11307), .Q(n6799) );
  NAND22 U2831 ( .A(n11329), .B(n11304), .Q(n6791) );
  NAND22 U2836 ( .A(n11329), .B(n11307), .Q(n6775) );
  NAND22 U2841 ( .A(n11325), .B(n11304), .Q(n6739) );
  NAND22 U2846 ( .A(n11325), .B(n11307), .Q(n6723) );
  NAND22 U2851 ( .A(n11338), .B(n11304), .Q(n6867) );
  NAND22 U2852 ( .A(n11338), .B(n11307), .Q(n6851) );
  NAND22 U2857 ( .A(n11324), .B(n11304), .Q(n6843) );
  NAND22 U2862 ( .A(n11324), .B(n11307), .Q(n6827) );
  NAND22 U2867 ( .A(n11333), .B(n11304), .Q(n6919) );
  NAND22 U2872 ( .A(n11333), .B(n11307), .Q(n6903) );
  NAND22 U2873 ( .A(n11328), .B(n11304), .Q(n6895) );
  NAND22 U2874 ( .A(n11328), .B(n11307), .Q(n6879) );
  NAND22 U2875 ( .A(n11336), .B(n11308), .Q(n6605) );
  NAND22 U2880 ( .A(n11336), .B(n11311), .Q(n6589) );
  NAND22 U2885 ( .A(n11331), .B(n11308), .Q(n6581) );
  NAND22 U2890 ( .A(n11331), .B(n11311), .Q(n6565) );
  NAND22 U2895 ( .A(n11337), .B(n11308), .Q(n6553) );
  NAND22 U2896 ( .A(n11337), .B(n11311), .Q(n6537) );
  NAND22 U2901 ( .A(n11327), .B(n11308), .Q(n6529) );
  NAND22 U2906 ( .A(n11327), .B(n11311), .Q(n6513) );
  NAND22 U2911 ( .A(n11340), .B(n11308), .Q(n6657) );
  NAND22 U2916 ( .A(n11340), .B(n11311), .Q(n6641) );
  NAND22 U2917 ( .A(n11326), .B(n11308), .Q(n6633) );
  NAND22 U2922 ( .A(n11326), .B(n11311), .Q(n6617) );
  NAND22 U2927 ( .A(n11335), .B(n11308), .Q(n6709) );
  NAND22 U2932 ( .A(n11335), .B(n11311), .Q(n6693) );
  NAND22 U2937 ( .A(n11334), .B(n11308), .Q(n6817) );
  NAND22 U2938 ( .A(n11334), .B(n11311), .Q(n6801) );
  NAND22 U2943 ( .A(n11329), .B(n11308), .Q(n6793) );
  NAND22 U2948 ( .A(n11329), .B(n11311), .Q(n6777) );
  NAND22 U2953 ( .A(n11325), .B(n11308), .Q(n6741) );
  NAND22 U2958 ( .A(n11325), .B(n11311), .Q(n6725) );
  NAND22 U2959 ( .A(n11338), .B(n11308), .Q(n6869) );
  NAND22 U2960 ( .A(n11338), .B(n11311), .Q(n6853) );
  NAND22 U2965 ( .A(n11324), .B(n11308), .Q(n6845) );
  NAND22 U2970 ( .A(n11324), .B(n11311), .Q(n6829) );
  NAND22 U2975 ( .A(n11333), .B(n11308), .Q(n6921) );
  NAND22 U2980 ( .A(n11333), .B(n11311), .Q(n6905) );
  NAND22 U2981 ( .A(n11328), .B(n11308), .Q(n6897) );
  NAND22 U2986 ( .A(n11328), .B(n11311), .Q(n6881) );
  NAND22 U2991 ( .A(n11336), .B(n11306), .Q(n6591) );
  NAND22 U2996 ( .A(n11331), .B(n11306), .Q(n6567) );
  NAND22 U3001 ( .A(n11337), .B(n11306), .Q(n6539) );
  NAND22 U3002 ( .A(n11327), .B(n11306), .Q(n6515) );
  NAND22 U3007 ( .A(n11340), .B(n11306), .Q(n6643) );
  NAND22 U3012 ( .A(n11326), .B(n11306), .Q(n6619) );
  NAND22 U3017 ( .A(n11335), .B(n11306), .Q(n6695) );
  NAND22 U3022 ( .A(n11334), .B(n11306), .Q(n6803) );
  NAND22 U3023 ( .A(n11329), .B(n11306), .Q(n6779) );
  NAND22 U3028 ( .A(n11325), .B(n11306), .Q(n6727) );
  NAND22 U3033 ( .A(n11338), .B(n11306), .Q(n6855) );
  NAND22 U3038 ( .A(n11324), .B(n11306), .Q(n6831) );
  NAND22 U3043 ( .A(n11333), .B(n11306), .Q(n6907) );
  NAND22 U3044 ( .A(n11328), .B(n11306), .Q(n6883) );
  NAND22 U3045 ( .A(n11309), .B(n11339), .Q(n6761) );
  NAND22 U3046 ( .A(n11305), .B(n11339), .Q(n6759) );
  NAND22 U3051 ( .A(n11304), .B(n11339), .Q(n6763) );
  NAND22 U3056 ( .A(n11308), .B(n11339), .Q(n6765) );
  NAND22 U3061 ( .A(n11311), .B(n11339), .Q(n6749) );
  NAND22 U3066 ( .A(n11307), .B(n11339), .Q(n6747) );
  NAND22 U3067 ( .A(n11306), .B(n11339), .Q(n6751) );
  NAND22 U3072 ( .A(n6146), .B(n11339), .Q(n6753) );
  NAND22 U3077 ( .A(n11309), .B(n11330), .Q(n6681) );
  NAND22 U3082 ( .A(n11305), .B(n11330), .Q(n6679) );
  NAND22 U3087 ( .A(n11304), .B(n11330), .Q(n6683) );
  NAND22 U3088 ( .A(n11308), .B(n11330), .Q(n6685) );
  NAND22 U3093 ( .A(n11311), .B(n11330), .Q(n6669) );
  NAND22 U3098 ( .A(n11307), .B(n11330), .Q(n6667) );
  NAND22 U3103 ( .A(n11306), .B(n11330), .Q(n6671) );
  INV3 U3108 ( .A(n10866), .Q(n11310) );
  NAND22 U3109 ( .A(n10857), .B(n10860), .Q(n10866) );
  NAND22 U3114 ( .A(n11336), .B(n6146), .Q(n6593) );
  NAND22 U3119 ( .A(n11337), .B(n6146), .Q(n6541) );
  NAND22 U3124 ( .A(n11340), .B(n6146), .Q(n6645) );
  NAND22 U3129 ( .A(n11335), .B(n6146), .Q(n6697) );
  NAND22 U3130 ( .A(n11329), .B(n6146), .Q(n6781) );
  NAND22 U3131 ( .A(n11331), .B(n6147), .Q(n6569) );
  NAND22 U3136 ( .A(n11327), .B(n6147), .Q(n6517) );
  NAND22 U3141 ( .A(n11326), .B(n6147), .Q(n6621) );
  NAND22 U3146 ( .A(n11334), .B(n6145), .Q(n6805) );
  NAND22 U3151 ( .A(n11325), .B(n6147), .Q(n6729) );
  NAND22 U3152 ( .A(n11338), .B(n6145), .Q(n6857) );
  NAND22 U3157 ( .A(n11324), .B(n6145), .Q(n6833) );
  NAND22 U3162 ( .A(n11333), .B(n6145), .Q(n6909) );
  NAND22 U3167 ( .A(n11328), .B(n6145), .Q(n6885) );
  NOR21 U3172 ( .A(n11347), .B(n11346), .Q(n6476) );
  NOR21 U3173 ( .A(n11345), .B(n11344), .Q(n6478) );
  NOR21 U3178 ( .A(n11351), .B(n11350), .Q(n6381) );
  NOR21 U3183 ( .A(n11349), .B(n11348), .Q(n6294) );
  NAND22 U3188 ( .A(n6480), .B(n6481), .Q(n6203) );
  NAND22 U3193 ( .A(n6487), .B(n6481), .Q(n6211) );
  NAND22 U3194 ( .A(n6493), .B(n6481), .Q(n6219) );
  NAND22 U3199 ( .A(n6480), .B(n6483), .Q(n6205) );
  NAND22 U3204 ( .A(n6487), .B(n6483), .Q(n6213) );
  NAND22 U3209 ( .A(n6493), .B(n6483), .Q(n6221) );
  NAND22 U3214 ( .A(n6476), .B(n6483), .Q(n6231) );
  NAND22 U3215 ( .A(n6480), .B(n6475), .Q(n6207) );
  NAND22 U3216 ( .A(n6487), .B(n6475), .Q(n6215) );
  NAND22 U3217 ( .A(n6481), .B(n6476), .Q(n6229) );
  NAND22 U3222 ( .A(n6475), .B(n6476), .Q(n6196) );
  NAND22 U3227 ( .A(n6480), .B(n6478), .Q(n6209) );
  NAND22 U3232 ( .A(n6487), .B(n6478), .Q(n6217) );
  NAND22 U3237 ( .A(n6475), .B(n6493), .Q(n6225) );
  NAND22 U3238 ( .A(n6478), .B(n6493), .Q(n6227) );
  NAND22 U3243 ( .A(n10860), .B(n10864), .Q(n10875) );
  NAND22 U3248 ( .A(n10855), .B(n10864), .Q(n10872) );
  NAND22 U3253 ( .A(n10855), .B(n10857), .Q(n10862) );
  NAND22 U3258 ( .A(n10874), .B(n10855), .Q(n10877) );
  NAND22 U3259 ( .A(n10874), .B(n10860), .Q(n10879) );
  NAND22 U3264 ( .A(n10852), .B(n10860), .Q(n10859) );
  NAND22 U3269 ( .A(n10852), .B(n10855), .Q(n10854) );
  NAND22 U3274 ( .A(n10783), .B(n10739), .Q(n10788) );
  NAND41 U3279 ( .A(n6555), .B(n6556), .C(n6557), .D(n6558), .Q(n6501) );
  NOR40 U3280 ( .A(n6559), .B(n6560), .C(n6561), .D(n6562), .Q(n6558) );
  NOR40 U3285 ( .A(n6571), .B(n6572), .C(n6573), .D(n6574), .Q(n6557) );
  NOR40 U3290 ( .A(n6583), .B(n6584), .C(n6585), .D(n6586), .Q(n6556) );
  NAND41 U3295 ( .A(n6767), .B(n6768), .C(n6769), .D(n6770), .Q(n6713) );
  NOR40 U3300 ( .A(n6771), .B(n6772), .C(n6773), .D(n6774), .Q(n6770) );
  NOR40 U3301 ( .A(n6783), .B(n6784), .C(n6785), .D(n6786), .Q(n6769) );
  NOR40 U3302 ( .A(n6795), .B(n6796), .C(n6797), .D(n6798), .Q(n6768) );
  NAND41 U3307 ( .A(n6949), .B(n6950), .C(n6951), .D(n6952), .Q(n6927) );
  NOR40 U3312 ( .A(n6953), .B(n6954), .C(n6955), .D(n6956), .Q(n6952) );
  NOR40 U3317 ( .A(n6957), .B(n6958), .C(n6959), .D(n6960), .Q(n6951) );
  NOR40 U3322 ( .A(n6961), .B(n6962), .C(n6963), .D(n6964), .Q(n6950) );
  NAND41 U3323 ( .A(n7033), .B(n7034), .C(n7035), .D(n7036), .Q(n7011) );
  NOR40 U3328 ( .A(n7037), .B(n7038), .C(n7039), .D(n7040), .Q(n7036) );
  NOR40 U3333 ( .A(n7041), .B(n7042), .C(n7043), .D(n7044), .Q(n7035) );
  NOR40 U3338 ( .A(n7045), .B(n7046), .C(n7047), .D(n7048), .Q(n7034) );
  NAND41 U3343 ( .A(n7119), .B(n7120), .C(n7121), .D(n7122), .Q(n7097) );
  NOR40 U3344 ( .A(n7123), .B(n7124), .C(n7125), .D(n7126), .Q(n7122) );
  NOR40 U3349 ( .A(n7127), .B(n7128), .C(n7129), .D(n7130), .Q(n7121) );
  NOR40 U3354 ( .A(n7131), .B(n7132), .C(n7133), .D(n7134), .Q(n7120) );
  NAND41 U3359 ( .A(n7203), .B(n7204), .C(n7205), .D(n7206), .Q(n7181) );
  NOR40 U3364 ( .A(n7207), .B(n7208), .C(n7209), .D(n7210), .Q(n7206) );
  NOR40 U3365 ( .A(n7211), .B(n7212), .C(n7213), .D(n7214), .Q(n7205) );
  NOR40 U3370 ( .A(n7215), .B(n7216), .C(n7217), .D(n7218), .Q(n7204) );
  NAND41 U3375 ( .A(n7289), .B(n7290), .C(n7291), .D(n7292), .Q(n7267) );
  NOR40 U3380 ( .A(n7293), .B(n7294), .C(n7295), .D(n7296), .Q(n7292) );
  NOR40 U3385 ( .A(n7297), .B(n7298), .C(n7299), .D(n7300), .Q(n7291) );
  NOR40 U3386 ( .A(n7301), .B(n7302), .C(n7303), .D(n7304), .Q(n7290) );
  NAND41 U3387 ( .A(n7373), .B(n7374), .C(n7375), .D(n7376), .Q(n7351) );
  NOR40 U3388 ( .A(n7377), .B(n7378), .C(n7379), .D(n7380), .Q(n7376) );
  NOR40 U3393 ( .A(n7381), .B(n7382), .C(n7383), .D(n7384), .Q(n7375) );
  NOR40 U3398 ( .A(n7385), .B(n7386), .C(n7387), .D(n7388), .Q(n7374) );
  NAND41 U3403 ( .A(n7459), .B(n7460), .C(n7461), .D(n7462), .Q(n7437) );
  NOR40 U3408 ( .A(n7463), .B(n7464), .C(n7465), .D(n7466), .Q(n7462) );
  NOR40 U3409 ( .A(n7467), .B(n7468), .C(n7469), .D(n7470), .Q(n7461) );
  NOR40 U3414 ( .A(n7471), .B(n7472), .C(n7473), .D(n7474), .Q(n7460) );
  NAND41 U3419 ( .A(n7543), .B(n7544), .C(n7545), .D(n7546), .Q(n7521) );
  NOR40 U3424 ( .A(n7547), .B(n7548), .C(n7549), .D(n7550), .Q(n7546) );
  NOR40 U3429 ( .A(n7551), .B(n7552), .C(n7553), .D(n7554), .Q(n7545) );
  NOR40 U3430 ( .A(n7555), .B(n7556), .C(n7557), .D(n7558), .Q(n7544) );
  NAND41 U3435 ( .A(n7629), .B(n7630), .C(n7631), .D(n7632), .Q(n7607) );
  NOR40 U3440 ( .A(n7633), .B(n7634), .C(n7635), .D(n7636), .Q(n7632) );
  NOR40 U3445 ( .A(n7637), .B(n7638), .C(n7639), .D(n7640), .Q(n7631) );
  NOR40 U3450 ( .A(n7641), .B(n7642), .C(n7643), .D(n7644), .Q(n7630) );
  NAND41 U3451 ( .A(n7713), .B(n7714), .C(n7715), .D(n7716), .Q(n7691) );
  NOR40 U3456 ( .A(n7717), .B(n7718), .C(n7719), .D(n7720), .Q(n7716) );
  NOR40 U3461 ( .A(n7721), .B(n7722), .C(n7723), .D(n7724), .Q(n7715) );
  NOR40 U3466 ( .A(n7725), .B(n7726), .C(n7727), .D(n7728), .Q(n7714) );
  NAND41 U3471 ( .A(n7799), .B(n7800), .C(n7801), .D(n7802), .Q(n7777) );
  NOR40 U3472 ( .A(n7803), .B(n7804), .C(n7805), .D(n7806), .Q(n7802) );
  NOR40 U3473 ( .A(n7807), .B(n7808), .C(n7809), .D(n7810), .Q(n7801) );
  NOR40 U3478 ( .A(n7811), .B(n7812), .C(n7813), .D(n7814), .Q(n7800) );
  NAND41 U3483 ( .A(n7883), .B(n7884), .C(n7885), .D(n7886), .Q(n7861) );
  NOR40 U3488 ( .A(n7887), .B(n7888), .C(n7889), .D(n7890), .Q(n7886) );
  NOR40 U3493 ( .A(n7891), .B(n7892), .C(n7893), .D(n7894), .Q(n7885) );
  NOR40 U3494 ( .A(n7895), .B(n7896), .C(n7897), .D(n7898), .Q(n7884) );
  NAND41 U3499 ( .A(n7969), .B(n7970), .C(n7971), .D(n7972), .Q(n7947) );
  NOR40 U3504 ( .A(n7973), .B(n7974), .C(n7975), .D(n7976), .Q(n7972) );
  NOR40 U3509 ( .A(n7977), .B(n7978), .C(n7979), .D(n7980), .Q(n7971) );
  NOR40 U3514 ( .A(n7981), .B(n7982), .C(n7983), .D(n7984), .Q(n7970) );
  NAND41 U3515 ( .A(n8053), .B(n8054), .C(n8055), .D(n8056), .Q(n8031) );
  NOR40 U3520 ( .A(n8057), .B(n8058), .C(n8059), .D(n8060), .Q(n8056) );
  NOR40 U3525 ( .A(n8061), .B(n8062), .C(n8063), .D(n8064), .Q(n8055) );
  NOR40 U3530 ( .A(n8065), .B(n8066), .C(n8067), .D(n8068), .Q(n8054) );
  NAND41 U3535 ( .A(n8139), .B(n8140), .C(n8141), .D(n8142), .Q(n8117) );
  NOR40 U3536 ( .A(n8143), .B(n8144), .C(n8145), .D(n8146), .Q(n8142) );
  NOR40 U3541 ( .A(n8147), .B(n8148), .C(n8149), .D(n8150), .Q(n8141) );
  NOR40 U3546 ( .A(n8151), .B(n8152), .C(n8153), .D(n8154), .Q(n8140) );
  NAND41 U3551 ( .A(n8223), .B(n8224), .C(n8225), .D(n8226), .Q(n8201) );
  NOR40 U3556 ( .A(n8227), .B(n8228), .C(n8229), .D(n8230), .Q(n8226) );
  NOR40 U3557 ( .A(n8231), .B(n8232), .C(n8233), .D(n8234), .Q(n8225) );
  NOR40 U3558 ( .A(n8235), .B(n8236), .C(n8237), .D(n8238), .Q(n8224) );
  NAND41 U3559 ( .A(n8309), .B(n8310), .C(n8311), .D(n8312), .Q(n8287) );
  NOR40 U3564 ( .A(n8313), .B(n8314), .C(n8315), .D(n8316), .Q(n8312) );
  NOR40 U3569 ( .A(n8317), .B(n8318), .C(n8319), .D(n8320), .Q(n8311) );
  NOR40 U3574 ( .A(n8321), .B(n8322), .C(n8323), .D(n8324), .Q(n8310) );
  NAND41 U3579 ( .A(n8393), .B(n8394), .C(n8395), .D(n8396), .Q(n8371) );
  NOR40 U3580 ( .A(n8397), .B(n8398), .C(n8399), .D(n8400), .Q(n8396) );
  NOR40 U3585 ( .A(n8401), .B(n8402), .C(n8403), .D(n8404), .Q(n8395) );
  NOR40 U3590 ( .A(n8405), .B(n8406), .C(n8407), .D(n8408), .Q(n8394) );
  NAND41 U3595 ( .A(n8479), .B(n8480), .C(n8481), .D(n8482), .Q(n8457) );
  NOR40 U3600 ( .A(n8483), .B(n8484), .C(n8485), .D(n8486), .Q(n8482) );
  NOR40 U3601 ( .A(n8487), .B(n8488), .C(n8489), .D(n8490), .Q(n8481) );
  NOR40 U3606 ( .A(n8491), .B(n8492), .C(n8493), .D(n8494), .Q(n8480) );
  NAND41 U3611 ( .A(n8563), .B(n8564), .C(n8565), .D(n8566), .Q(n8541) );
  NOR40 U3616 ( .A(n8567), .B(n8568), .C(n8569), .D(n8570), .Q(n8566) );
  NOR40 U3621 ( .A(n8571), .B(n8572), .C(n8573), .D(n8574), .Q(n8565) );
  NOR40 U3622 ( .A(n8575), .B(n8576), .C(n8577), .D(n8578), .Q(n8564) );
  NAND41 U3627 ( .A(n8649), .B(n8650), .C(n8651), .D(n8652), .Q(n8627) );
  NOR40 U3632 ( .A(n8653), .B(n8654), .C(n8655), .D(n8656), .Q(n8652) );
  NOR40 U3637 ( .A(n8657), .B(n8658), .C(n8659), .D(n8660), .Q(n8651) );
  NOR40 U3642 ( .A(n8661), .B(n8662), .C(n8663), .D(n8664), .Q(n8650) );
  NAND41 U3643 ( .A(n8733), .B(n8734), .C(n8735), .D(n8736), .Q(n8711) );
  NOR40 U3644 ( .A(n8737), .B(n8738), .C(n8739), .D(n8740), .Q(n8736) );
  NOR40 U3649 ( .A(n8741), .B(n8742), .C(n8743), .D(n8744), .Q(n8735) );
  NOR40 U3654 ( .A(n8745), .B(n8746), .C(n8747), .D(n8748), .Q(n8734) );
  NAND41 U3659 ( .A(n8819), .B(n8820), .C(n8821), .D(n8822), .Q(n8797) );
  NOR40 U3664 ( .A(n8823), .B(n8824), .C(n8825), .D(n8826), .Q(n8822) );
  NOR40 U3665 ( .A(n8827), .B(n8828), .C(n8829), .D(n8830), .Q(n8821) );
  NOR40 U3670 ( .A(n8831), .B(n8832), .C(n8833), .D(n8834), .Q(n8820) );
  NAND41 U3675 ( .A(n8903), .B(n8904), .C(n8905), .D(n8906), .Q(n8881) );
  NOR40 U3680 ( .A(n8907), .B(n8908), .C(n8909), .D(n8910), .Q(n8906) );
  NOR40 U3685 ( .A(n8911), .B(n8912), .C(n8913), .D(n8914), .Q(n8905) );
  NOR40 U3686 ( .A(n8915), .B(n8916), .C(n8917), .D(n8918), .Q(n8904) );
  NAND41 U3691 ( .A(n8989), .B(n8990), .C(n8991), .D(n8992), .Q(n8967) );
  NOR40 U3696 ( .A(n8993), .B(n8994), .C(n8995), .D(n8996), .Q(n8992) );
  NOR40 U3701 ( .A(n8997), .B(n8998), .C(n8999), .D(n9000), .Q(n8991) );
  NOR40 U3706 ( .A(n9001), .B(n9002), .C(n9003), .D(n9004), .Q(n8990) );
  NAND41 U3707 ( .A(n9073), .B(n9074), .C(n9075), .D(n9076), .Q(n9051) );
  NOR40 U3712 ( .A(n9077), .B(n9078), .C(n9079), .D(n9080), .Q(n9076) );
  NOR40 U3717 ( .A(n9081), .B(n9082), .C(n9083), .D(n9084), .Q(n9075) );
  NOR40 U3722 ( .A(n9085), .B(n9086), .C(n9087), .D(n9088), .Q(n9074) );
  NAND41 U3727 ( .A(n9159), .B(n9160), .C(n9161), .D(n9162), .Q(n9137) );
  NOR40 U3728 ( .A(n9163), .B(n9164), .C(n9165), .D(n9166), .Q(n9162) );
  NOR40 U3729 ( .A(n9167), .B(n9168), .C(n9169), .D(n9170), .Q(n9161) );
  NOR40 U3730 ( .A(n9171), .B(n9172), .C(n9173), .D(n9174), .Q(n9160) );
  NAND41 U3735 ( .A(n9243), .B(n9244), .C(n9245), .D(n9246), .Q(n9221) );
  NOR40 U3740 ( .A(n9247), .B(n9248), .C(n9249), .D(n9250), .Q(n9246) );
  NOR40 U3745 ( .A(n9251), .B(n9252), .C(n9253), .D(n9254), .Q(n9245) );
  NOR40 U3750 ( .A(n9255), .B(n9256), .C(n9257), .D(n9258), .Q(n9244) );
  NAND41 U3751 ( .A(n9329), .B(n9330), .C(n9331), .D(n9332), .Q(n9307) );
  NOR40 U3756 ( .A(n9333), .B(n9334), .C(n9335), .D(n9336), .Q(n9332) );
  NOR40 U3761 ( .A(n9337), .B(n9338), .C(n9339), .D(n9340), .Q(n9331) );
  NOR40 U3766 ( .A(n9341), .B(n9342), .C(n9343), .D(n9344), .Q(n9330) );
  NAND41 U3771 ( .A(n9413), .B(n9414), .C(n9415), .D(n9416), .Q(n9391) );
  NOR40 U3772 ( .A(n9417), .B(n9418), .C(n9419), .D(n9420), .Q(n9416) );
  NOR40 U3777 ( .A(n9421), .B(n9422), .C(n9423), .D(n9424), .Q(n9415) );
  NOR40 U3782 ( .A(n9425), .B(n9426), .C(n9427), .D(n9428), .Q(n9414) );
  NAND41 U3787 ( .A(n9499), .B(n9500), .C(n9501), .D(n9502), .Q(n9477) );
  NOR40 U3792 ( .A(n9503), .B(n9504), .C(n9505), .D(n9506), .Q(n9502) );
  NOR40 U3793 ( .A(n9507), .B(n9508), .C(n9509), .D(n9510), .Q(n9501) );
  NOR40 U3798 ( .A(n9511), .B(n9512), .C(n9513), .D(n9514), .Q(n9500) );
  NAND41 U3803 ( .A(n9583), .B(n9584), .C(n9585), .D(n9586), .Q(n9561) );
  NOR40 U3808 ( .A(n9587), .B(n9588), .C(n9589), .D(n9590), .Q(n9586) );
  NOR40 U3813 ( .A(n9591), .B(n9592), .C(n9593), .D(n9594), .Q(n9585) );
  NOR40 U3814 ( .A(n9595), .B(n9596), .C(n9597), .D(n9598), .Q(n9584) );
  NAND41 U3815 ( .A(n9669), .B(n9670), .C(n9671), .D(n9672), .Q(n9647) );
  NOR40 U3820 ( .A(n9673), .B(n9674), .C(n9675), .D(n9676), .Q(n9672) );
  NOR40 U3825 ( .A(n9677), .B(n9678), .C(n9679), .D(n9680), .Q(n9671) );
  NOR40 U3830 ( .A(n9681), .B(n9682), .C(n9683), .D(n9684), .Q(n9670) );
  NAND41 U3835 ( .A(n9753), .B(n9754), .C(n9755), .D(n9756), .Q(n9731) );
  NOR40 U3836 ( .A(n9757), .B(n9758), .C(n9759), .D(n9760), .Q(n9756) );
  NOR40 U3841 ( .A(n9761), .B(n9762), .C(n9763), .D(n9764), .Q(n9755) );
  NOR40 U3846 ( .A(n9765), .B(n9766), .C(n9767), .D(n9768), .Q(n9754) );
  NAND41 U3851 ( .A(n9839), .B(n9840), .C(n9841), .D(n9842), .Q(n9817) );
  NOR40 U3856 ( .A(n9843), .B(n9844), .C(n9845), .D(n9846), .Q(n9842) );
  NOR40 U3857 ( .A(n9847), .B(n9848), .C(n9849), .D(n9850), .Q(n9841) );
  NOR40 U3862 ( .A(n9851), .B(n9852), .C(n9853), .D(n9854), .Q(n9840) );
  NAND41 U3867 ( .A(n9923), .B(n9924), .C(n9925), .D(n9926), .Q(n9901) );
  NOR40 U3872 ( .A(n9927), .B(n9928), .C(n9929), .D(n9930), .Q(n9926) );
  NOR40 U3877 ( .A(n9931), .B(n9932), .C(n9933), .D(n9934), .Q(n9925) );
  NOR40 U3878 ( .A(n9935), .B(n9936), .C(n9937), .D(n9938), .Q(n9924) );
  NAND41 U3883 ( .A(n10009), .B(n10010), .C(n10011), .D(n10012), .Q(n9987) );
  NOR40 U3888 ( .A(n10013), .B(n10014), .C(n10015), .D(n10016), .Q(n10012) );
  NOR40 U3893 ( .A(n10017), .B(n10018), .C(n10019), .D(n10020), .Q(n10011) );
  NOR40 U3898 ( .A(n10021), .B(n10022), .C(n10023), .D(n10024), .Q(n10010) );
  NAND41 U3899 ( .A(n10093), .B(n10094), .C(n10095), .D(n10096), .Q(n10071) );
  NOR40 U3900 ( .A(n10097), .B(n10098), .C(n10099), .D(n10100), .Q(n10096) );
  NOR40 U3901 ( .A(n10101), .B(n10102), .C(n10103), .D(n10104), .Q(n10095) );
  NOR40 U3906 ( .A(n10105), .B(n10106), .C(n10107), .D(n10108), .Q(n10094) );
  NAND41 U3911 ( .A(n10179), .B(n10180), .C(n10181), .D(n10182), .Q(n10157) );
  NOR40 U3916 ( .A(n10183), .B(n10184), .C(n10185), .D(n10186), .Q(n10182) );
  NOR40 U3921 ( .A(n10187), .B(n10188), .C(n10189), .D(n10190), .Q(n10181) );
  NOR40 U3922 ( .A(n10191), .B(n10192), .C(n10193), .D(n10194), .Q(n10180) );
  NAND41 U3927 ( .A(n10263), .B(n10264), .C(n10265), .D(n10266), .Q(n10241) );
  NOR40 U3932 ( .A(n10267), .B(n10268), .C(n10269), .D(n10270), .Q(n10266) );
  NOR40 U3937 ( .A(n10271), .B(n10272), .C(n10273), .D(n10274), .Q(n10265) );
  NOR40 U3942 ( .A(n10275), .B(n10276), .C(n10277), .D(n10278), .Q(n10264) );
  NAND41 U3943 ( .A(n10349), .B(n10350), .C(n10351), .D(n10352), .Q(n10327) );
  NOR40 U3948 ( .A(n10353), .B(n10354), .C(n10355), .D(n10356), .Q(n10352) );
  NOR40 U3953 ( .A(n10357), .B(n10358), .C(n10359), .D(n10360), .Q(n10351) );
  NOR40 U3958 ( .A(n10361), .B(n10362), .C(n10363), .D(n10364), .Q(n10350) );
  NAND41 U3963 ( .A(n10433), .B(n10434), .C(n10435), .D(n10436), .Q(n10411) );
  NOR40 U3964 ( .A(n10437), .B(n10438), .C(n10439), .D(n10440), .Q(n10436) );
  NOR40 U3969 ( .A(n10441), .B(n10442), .C(n10443), .D(n10444), .Q(n10435) );
  NOR40 U3974 ( .A(n10445), .B(n10446), .C(n10447), .D(n10448), .Q(n10434) );
  NAND41 U3979 ( .A(n10519), .B(n10520), .C(n10521), .D(n10522), .Q(n10497) );
  NOR40 U3984 ( .A(n10523), .B(n10524), .C(n10525), .D(n10526), .Q(n10522) );
  NOR40 U3985 ( .A(n10527), .B(n10528), .C(n10529), .D(n10530), .Q(n10521) );
  NOR40 U3986 ( .A(n10531), .B(n10532), .C(n10533), .D(n10534), .Q(n10520) );
  NAND41 U3991 ( .A(n10603), .B(n10604), .C(n10605), .D(n10606), .Q(n10581) );
  NOR40 U3996 ( .A(n10607), .B(n10608), .C(n10609), .D(n10610), .Q(n10606) );
  NOR40 U4001 ( .A(n10611), .B(n10612), .C(n10613), .D(n10614), .Q(n10605) );
  NOR40 U4006 ( .A(n10615), .B(n10616), .C(n10617), .D(n10618), .Q(n10604) );
  NAND41 U4007 ( .A(n10692), .B(n10693), .C(n10694), .D(n10695), .Q(n10667) );
  NOR40 U4012 ( .A(n10696), .B(n10697), .C(n10698), .D(n10699), .Q(n10695) );
  NOR40 U4017 ( .A(n10700), .B(n10701), .C(n10702), .D(n10703), .Q(n10694) );
  NOR40 U4022 ( .A(n10704), .B(n10705), .C(n10706), .D(n10707), .Q(n10693) );
  NAND41 U4027 ( .A(n10789), .B(n10790), .C(n10791), .D(n10792), .Q(n10764) );
  NOR40 U4028 ( .A(n10793), .B(n10794), .C(n10795), .D(n10796), .Q(n10792) );
  NOR40 U4033 ( .A(n10797), .B(n10798), .C(n10799), .D(n10800), .Q(n10791) );
  NOR40 U4038 ( .A(n10801), .B(n10802), .C(n10803), .D(n10804), .Q(n10790) );
  NAND41 U4043 ( .A(n6503), .B(n6504), .C(n6505), .D(n6506), .Q(n6502) );
  NOR40 U4048 ( .A(n6507), .B(n6508), .C(n6509), .D(n6510), .Q(n6506) );
  NOR40 U4049 ( .A(n6519), .B(n6520), .C(n6521), .D(n6522), .Q(n6505) );
  NOR40 U4054 ( .A(n6531), .B(n6532), .C(n6533), .D(n6534), .Q(n6504) );
  NAND41 U4059 ( .A(n6607), .B(n6608), .C(n6609), .D(n6610), .Q(n6500) );
  NOR40 U4064 ( .A(n6611), .B(n6612), .C(n6613), .D(n6614), .Q(n6610) );
  NOR40 U4069 ( .A(n6623), .B(n6624), .C(n6625), .D(n6626), .Q(n6609) );
  NOR40 U4070 ( .A(n6635), .B(n6636), .C(n6637), .D(n6638), .Q(n6608) );
  NAND41 U4071 ( .A(n6715), .B(n6716), .C(n6717), .D(n6718), .Q(n6714) );
  NOR40 U4072 ( .A(n6719), .B(n6720), .C(n6721), .D(n6722), .Q(n6718) );
  NOR40 U4077 ( .A(n6731), .B(n6732), .C(n6733), .D(n6734), .Q(n6717) );
  NOR40 U4082 ( .A(n6743), .B(n6744), .C(n6745), .D(n6746), .Q(n6716) );
  NAND41 U4087 ( .A(n6819), .B(n6820), .C(n6821), .D(n6822), .Q(n6712) );
  NOR40 U4092 ( .A(n6823), .B(n6824), .C(n6825), .D(n6826), .Q(n6822) );
  NOR40 U4093 ( .A(n6835), .B(n6836), .C(n6837), .D(n6838), .Q(n6821) );
  NOR40 U4098 ( .A(n6847), .B(n6848), .C(n6849), .D(n6850), .Q(n6820) );
  NAND41 U4103 ( .A(n6929), .B(n6930), .C(n6931), .D(n6932), .Q(n6928) );
  NOR40 U4108 ( .A(n6933), .B(n6934), .C(n6935), .D(n6936), .Q(n6932) );
  NOR40 U4113 ( .A(n6937), .B(n6938), .C(n6939), .D(n6940), .Q(n6931) );
  NOR40 U4114 ( .A(n6941), .B(n6942), .C(n6943), .D(n6944), .Q(n6930) );
  NAND41 U4119 ( .A(n6969), .B(n6970), .C(n6971), .D(n6972), .Q(n6926) );
  NOR40 U4124 ( .A(n6973), .B(n6974), .C(n6975), .D(n6976), .Q(n6972) );
  NOR40 U4129 ( .A(n6977), .B(n6978), .C(n6979), .D(n6980), .Q(n6971) );
  NOR40 U4134 ( .A(n6981), .B(n6982), .C(n6983), .D(n6984), .Q(n6970) );
  NAND41 U4135 ( .A(n7013), .B(n7014), .C(n7015), .D(n7016), .Q(n7012) );
  NOR40 U4140 ( .A(n7017), .B(n7018), .C(n7019), .D(n7020), .Q(n7016) );
  NOR40 U4145 ( .A(n7021), .B(n7022), .C(n7023), .D(n7024), .Q(n7015) );
  NOR40 U4150 ( .A(n7025), .B(n7026), .C(n7027), .D(n7028), .Q(n7014) );
  NAND41 U4155 ( .A(n7053), .B(n7054), .C(n7055), .D(n7056), .Q(n7010) );
  NOR40 U4156 ( .A(n7057), .B(n7058), .C(n7059), .D(n7060), .Q(n7056) );
  NOR40 U4157 ( .A(n7061), .B(n7062), .C(n7063), .D(n7064), .Q(n7055) );
  NOR40 U4162 ( .A(n7065), .B(n7066), .C(n7067), .D(n7068), .Q(n7054) );
  NAND41 U4167 ( .A(n7099), .B(n7100), .C(n7101), .D(n7102), .Q(n7098) );
  NOR40 U4172 ( .A(n7103), .B(n7104), .C(n7105), .D(n7106), .Q(n7102) );
  NOR40 U4177 ( .A(n7107), .B(n7108), .C(n7109), .D(n7110), .Q(n7101) );
  NOR40 U4178 ( .A(n7111), .B(n7112), .C(n7113), .D(n7114), .Q(n7100) );
  NAND41 U4183 ( .A(n7139), .B(n7140), .C(n7141), .D(n7142), .Q(n7096) );
  NOR40 U4188 ( .A(n7143), .B(n7144), .C(n7145), .D(n7146), .Q(n7142) );
  NOR40 U4193 ( .A(n7147), .B(n7148), .C(n7149), .D(n7150), .Q(n7141) );
  NOR40 U4198 ( .A(n7151), .B(n7152), .C(n7153), .D(n7154), .Q(n7140) );
  NAND41 U4199 ( .A(n7183), .B(n7184), .C(n7185), .D(n7186), .Q(n7182) );
  NOR40 U4204 ( .A(n7187), .B(n7188), .C(n7189), .D(n7190), .Q(n7186) );
  NOR40 U4209 ( .A(n7191), .B(n7192), .C(n7193), .D(n7194), .Q(n7185) );
  NOR40 U4214 ( .A(n7195), .B(n7196), .C(n7197), .D(n7198), .Q(n7184) );
  NAND41 U4219 ( .A(n7223), .B(n7224), .C(n7225), .D(n7226), .Q(n7180) );
  NOR40 U4220 ( .A(n7227), .B(n7228), .C(n7229), .D(n7230), .Q(n7226) );
  NOR40 U4225 ( .A(n7231), .B(n7232), .C(n7233), .D(n7234), .Q(n7225) );
  NOR40 U4230 ( .A(n7235), .B(n7236), .C(n7237), .D(n7238), .Q(n7224) );
  NAND41 U4235 ( .A(n7269), .B(n7270), .C(n7271), .D(n7272), .Q(n7268) );
  NOR40 U4240 ( .A(n7273), .B(n7274), .C(n7275), .D(n7276), .Q(n7272) );
  NOR40 U4241 ( .A(n7277), .B(n7278), .C(n7279), .D(n7280), .Q(n7271) );
  NOR40 U4242 ( .A(n7281), .B(n7282), .C(n7283), .D(n7284), .Q(n7270) );
  NAND41 U4243 ( .A(n7309), .B(n7310), .C(n7311), .D(n7312), .Q(n7266) );
  NOR40 U4245 ( .A(n7313), .B(n7314), .C(n7315), .D(n7316), .Q(n7312) );
  NOR40 U4246 ( .A(n7317), .B(n7318), .C(n7319), .D(n7320), .Q(n7311) );
  NOR40 U4248 ( .A(n7321), .B(n7322), .C(n7323), .D(n7324), .Q(n7310) );
  NAND41 U4249 ( .A(n7353), .B(n7354), .C(n7355), .D(n7356), .Q(n7352) );
  NOR40 U4251 ( .A(n7357), .B(n7358), .C(n7359), .D(n7360), .Q(n7356) );
  NOR40 U4252 ( .A(n7361), .B(n7362), .C(n7363), .D(n7364), .Q(n7355) );
  NOR40 U4254 ( .A(n7365), .B(n7366), .C(n7367), .D(n7368), .Q(n7354) );
  NAND41 U4255 ( .A(n7393), .B(n7394), .C(n7395), .D(n7396), .Q(n7350) );
  NOR40 U4256 ( .A(n7397), .B(n7398), .C(n7399), .D(n7400), .Q(n7396) );
  NOR40 U4258 ( .A(n7401), .B(n7402), .C(n7403), .D(n7404), .Q(n7395) );
  NOR40 U4259 ( .A(n7405), .B(n7406), .C(n7407), .D(n7408), .Q(n7394) );
  NAND41 U4261 ( .A(n7439), .B(n7440), .C(n7441), .D(n7442), .Q(n7438) );
  NOR40 U4262 ( .A(n7443), .B(n7444), .C(n7445), .D(n7446), .Q(n7442) );
  NOR40 U4264 ( .A(n7447), .B(n7448), .C(n7449), .D(n7450), .Q(n7441) );
  NOR40 U4265 ( .A(n7451), .B(n7452), .C(n7453), .D(n7454), .Q(n7440) );
  NAND41 U4267 ( .A(n7479), .B(n7480), .C(n7481), .D(n7482), .Q(n7436) );
  NOR40 U4268 ( .A(n7483), .B(n7484), .C(n7485), .D(n7486), .Q(n7482) );
  NOR40 U4269 ( .A(n7487), .B(n7488), .C(n7489), .D(n7490), .Q(n7481) );
  NOR40 U4271 ( .A(n7491), .B(n7492), .C(n7493), .D(n7494), .Q(n7480) );
  NAND41 U4272 ( .A(n7523), .B(n7524), .C(n7525), .D(n7526), .Q(n7522) );
  NOR40 U4274 ( .A(n7527), .B(n7528), .C(n7529), .D(n7530), .Q(n7526) );
  NOR40 U4275 ( .A(n7531), .B(n7532), .C(n7533), .D(n7534), .Q(n7525) );
  NOR40 U4277 ( .A(n7535), .B(n7536), .C(n7537), .D(n7538), .Q(n7524) );
  NAND41 U4278 ( .A(n7563), .B(n7564), .C(n7565), .D(n7566), .Q(n7520) );
  NOR40 U4280 ( .A(n7567), .B(n7568), .C(n7569), .D(n7570), .Q(n7566) );
  NOR40 U4281 ( .A(n7571), .B(n7572), .C(n7573), .D(n7574), .Q(n7565) );
  NOR40 U4282 ( .A(n7575), .B(n7576), .C(n7577), .D(n7578), .Q(n7564) );
  NAND41 U4283 ( .A(n7609), .B(n7610), .C(n7611), .D(n7612), .Q(n7608) );
  NOR40 U4285 ( .A(n7613), .B(n7614), .C(n7615), .D(n7616), .Q(n7612) );
  NOR40 U4286 ( .A(n7617), .B(n7618), .C(n7619), .D(n7620), .Q(n7611) );
  NOR40 U4288 ( .A(n7621), .B(n7622), .C(n7623), .D(n7624), .Q(n7610) );
  NAND41 U4289 ( .A(n7649), .B(n7650), .C(n7651), .D(n7652), .Q(n7606) );
  NOR40 U4291 ( .A(n7653), .B(n7654), .C(n7655), .D(n7656), .Q(n7652) );
  NOR40 U4292 ( .A(n7657), .B(n7658), .C(n7659), .D(n7660), .Q(n7651) );
  NOR40 U4294 ( .A(n7661), .B(n7662), .C(n7663), .D(n7664), .Q(n7650) );
  NAND41 U4295 ( .A(n7693), .B(n7694), .C(n7695), .D(n7696), .Q(n7692) );
  NOR40 U4296 ( .A(n7697), .B(n7698), .C(n7699), .D(n7700), .Q(n7696) );
  NOR40 U4297 ( .A(n7701), .B(n7702), .C(n7703), .D(n7704), .Q(n7695) );
  NOR40 U4299 ( .A(n7705), .B(n7706), .C(n7707), .D(n7708), .Q(n7694) );
  NAND41 U4300 ( .A(n7733), .B(n7734), .C(n7735), .D(n7736), .Q(n7690) );
  NOR40 U4302 ( .A(n7737), .B(n7738), .C(n7739), .D(n7740), .Q(n7736) );
  NOR40 U4303 ( .A(n7741), .B(n7742), .C(n7743), .D(n7744), .Q(n7735) );
  NOR40 U4305 ( .A(n7745), .B(n7746), .C(n7747), .D(n7748), .Q(n7734) );
  NAND41 U4306 ( .A(n7779), .B(n7780), .C(n7781), .D(n7782), .Q(n7778) );
  NOR40 U4308 ( .A(n7783), .B(n7784), .C(n7785), .D(n7786), .Q(n7782) );
  NOR40 U4309 ( .A(n7787), .B(n7788), .C(n7789), .D(n7790), .Q(n7781) );
  NOR40 U4310 ( .A(n7791), .B(n7792), .C(n7793), .D(n7794), .Q(n7780) );
  NAND41 U4312 ( .A(n7819), .B(n7820), .C(n7821), .D(n7822), .Q(n7776) );
  NOR40 U4313 ( .A(n7823), .B(n7824), .C(n7825), .D(n7826), .Q(n7822) );
  NOR40 U4315 ( .A(n7827), .B(n7828), .C(n7829), .D(n7830), .Q(n7821) );
  NOR40 U4316 ( .A(n7831), .B(n7832), .C(n7833), .D(n7834), .Q(n7820) );
  NAND41 U4318 ( .A(n7863), .B(n7864), .C(n7865), .D(n7866), .Q(n7862) );
  NOR40 U4319 ( .A(n7867), .B(n7868), .C(n7869), .D(n7870), .Q(n7866) );
  NOR40 U4321 ( .A(n7871), .B(n7872), .C(n7873), .D(n7874), .Q(n7865) );
  NOR40 U4322 ( .A(n7875), .B(n7876), .C(n7877), .D(n7878), .Q(n7864) );
  NAND41 U4323 ( .A(n7903), .B(n7904), .C(n7905), .D(n7906), .Q(n7860) );
  NOR40 U4325 ( .A(n7907), .B(n7908), .C(n7909), .D(n7910), .Q(n7906) );
  NOR40 U4326 ( .A(n7911), .B(n7912), .C(n7913), .D(n7914), .Q(n7905) );
  NOR40 U4328 ( .A(n7915), .B(n7916), .C(n7917), .D(n7918), .Q(n7904) );
  NAND41 U4329 ( .A(n7949), .B(n7950), .C(n7951), .D(n7952), .Q(n7948) );
  NOR40 U4331 ( .A(n7953), .B(n7954), .C(n7955), .D(n7956), .Q(n7952) );
  NOR40 U4332 ( .A(n7957), .B(n7958), .C(n7959), .D(n7960), .Q(n7951) );
  NOR40 U4334 ( .A(n7961), .B(n7962), .C(n7963), .D(n7964), .Q(n7950) );
  NAND41 U4335 ( .A(n7989), .B(n7990), .C(n7991), .D(n7992), .Q(n7946) );
  NOR40 U4336 ( .A(n7993), .B(n7994), .C(n7995), .D(n7996), .Q(n7992) );
  NOR40 U4337 ( .A(n7997), .B(n7998), .C(n7999), .D(n8000), .Q(n7991) );
  NOR40 U4339 ( .A(n8001), .B(n8002), .C(n8003), .D(n8004), .Q(n7990) );
  NAND41 U4340 ( .A(n8033), .B(n8034), .C(n8035), .D(n8036), .Q(n8032) );
  NOR40 U4342 ( .A(n8037), .B(n8038), .C(n8039), .D(n8040), .Q(n8036) );
  NOR40 U4343 ( .A(n8041), .B(n8042), .C(n8043), .D(n8044), .Q(n8035) );
  NOR40 U4345 ( .A(n8045), .B(n8046), .C(n8047), .D(n8048), .Q(n8034) );
  NAND41 U4346 ( .A(n8073), .B(n8074), .C(n8075), .D(n8076), .Q(n8030) );
  NOR40 U4348 ( .A(n8077), .B(n8078), .C(n8079), .D(n8080), .Q(n8076) );
  NOR40 U4349 ( .A(n8081), .B(n8082), .C(n8083), .D(n8084), .Q(n8075) );
  NOR40 U4350 ( .A(n8085), .B(n8086), .C(n8087), .D(n8088), .Q(n8074) );
  NAND41 U4351 ( .A(n8119), .B(n8120), .C(n8121), .D(n8122), .Q(n8118) );
  NOR40 U4352 ( .A(n8123), .B(n8124), .C(n8125), .D(n8126), .Q(n8122) );
  NOR40 U4354 ( .A(n8127), .B(n8128), .C(n8129), .D(n8130), .Q(n8121) );
  NOR40 U4355 ( .A(n8131), .B(n8132), .C(n8133), .D(n8134), .Q(n8120) );
  NAND41 U4357 ( .A(n8159), .B(n8160), .C(n8161), .D(n8162), .Q(n8116) );
  NOR40 U4358 ( .A(n8163), .B(n8164), .C(n8165), .D(n8166), .Q(n8162) );
  NOR40 U4360 ( .A(n8167), .B(n8168), .C(n8169), .D(n8170), .Q(n8161) );
  NOR40 U4361 ( .A(n8171), .B(n8172), .C(n8173), .D(n8174), .Q(n8160) );
  NAND41 U4363 ( .A(n8203), .B(n8204), .C(n8205), .D(n8206), .Q(n8202) );
  NOR40 U4364 ( .A(n8207), .B(n8208), .C(n8209), .D(n8210), .Q(n8206) );
  NOR40 U4365 ( .A(n8211), .B(n8212), .C(n8213), .D(n8214), .Q(n8205) );
  NOR40 U4367 ( .A(n8215), .B(n8216), .C(n8217), .D(n8218), .Q(n8204) );
  NAND41 U4368 ( .A(n8243), .B(n8244), .C(n8245), .D(n8246), .Q(n8200) );
  NOR40 U4370 ( .A(n8247), .B(n8248), .C(n8249), .D(n8250), .Q(n8246) );
  NOR40 U4371 ( .A(n8251), .B(n8252), .C(n8253), .D(n8254), .Q(n8245) );
  NOR40 U4373 ( .A(n8255), .B(n8256), .C(n8257), .D(n8258), .Q(n8244) );
  NAND41 U4374 ( .A(n8289), .B(n8290), .C(n8291), .D(n8292), .Q(n8288) );
  NOR40 U4376 ( .A(n8293), .B(n8294), .C(n8295), .D(n8296), .Q(n8292) );
  NOR40 U4377 ( .A(n8297), .B(n8298), .C(n8299), .D(n8300), .Q(n8291) );
  NOR40 U4378 ( .A(n8301), .B(n8302), .C(n8303), .D(n8304), .Q(n8290) );
  NAND41 U4380 ( .A(n8329), .B(n8330), .C(n8331), .D(n8332), .Q(n8286) );
  NOR40 U4381 ( .A(n8333), .B(n8334), .C(n8335), .D(n8336), .Q(n8332) );
  NOR40 U4383 ( .A(n8337), .B(n8338), .C(n8339), .D(n8340), .Q(n8331) );
  NOR40 U4384 ( .A(n8341), .B(n8342), .C(n8343), .D(n8344), .Q(n8330) );
  NAND41 U4386 ( .A(n8373), .B(n8374), .C(n8375), .D(n8376), .Q(n8372) );
  NOR40 U4387 ( .A(n8377), .B(n8378), .C(n8379), .D(n8380), .Q(n8376) );
  NOR40 U4389 ( .A(n8381), .B(n8382), .C(n8383), .D(n8384), .Q(n8375) );
  NOR40 U4390 ( .A(n8385), .B(n8386), .C(n8387), .D(n8388), .Q(n8374) );
  NAND41 U4391 ( .A(n8413), .B(n8414), .C(n8415), .D(n8416), .Q(n8370) );
  NOR40 U4392 ( .A(n8417), .B(n8418), .C(n8419), .D(n8420), .Q(n8416) );
  NOR40 U4394 ( .A(n8421), .B(n8422), .C(n8423), .D(n8424), .Q(n8415) );
  NOR40 U4395 ( .A(n8425), .B(n8426), .C(n8427), .D(n8428), .Q(n8414) );
  NAND41 U4397 ( .A(n8459), .B(n8460), .C(n8461), .D(n8462), .Q(n8458) );
  NOR40 U4398 ( .A(n8463), .B(n8464), .C(n8465), .D(n8466), .Q(n8462) );
  NOR40 U4400 ( .A(n8467), .B(n8468), .C(n8469), .D(n8470), .Q(n8461) );
  NOR40 U4401 ( .A(n8471), .B(n8472), .C(n8473), .D(n8474), .Q(n8460) );
  NAND41 U4403 ( .A(n8499), .B(n8500), .C(n8501), .D(n8502), .Q(n8456) );
  NOR40 U4404 ( .A(n8503), .B(n8504), .C(n8505), .D(n8506), .Q(n8502) );
  NOR40 U4405 ( .A(n8507), .B(n8508), .C(n8509), .D(n8510), .Q(n8501) );
  NOR40 U4406 ( .A(n8511), .B(n8512), .C(n8513), .D(n8514), .Q(n8500) );
  NAND41 U4407 ( .A(n8543), .B(n8544), .C(n8545), .D(n8546), .Q(n8542) );
  NOR40 U4409 ( .A(n8547), .B(n8548), .C(n8549), .D(n8550), .Q(n8546) );
  NOR40 U4410 ( .A(n8551), .B(n8552), .C(n8553), .D(n8554), .Q(n8545) );
  NOR40 U4412 ( .A(n8555), .B(n8556), .C(n8557), .D(n8558), .Q(n8544) );
  NAND41 U4413 ( .A(n8583), .B(n8584), .C(n8585), .D(n8586), .Q(n8540) );
  NOR40 U4415 ( .A(n8587), .B(n8588), .C(n8589), .D(n8590), .Q(n8586) );
  NOR40 U4416 ( .A(n8591), .B(n8592), .C(n8593), .D(n8594), .Q(n8585) );
  NOR40 U4418 ( .A(n8595), .B(n8596), .C(n8597), .D(n8598), .Q(n8584) );
  NAND41 U4419 ( .A(n8629), .B(n8630), .C(n8631), .D(n8632), .Q(n8628) );
  NOR40 U4420 ( .A(n8633), .B(n8634), .C(n8635), .D(n8636), .Q(n8632) );
  NOR40 U4422 ( .A(n8637), .B(n8638), .C(n8639), .D(n8640), .Q(n8631) );
  NOR40 U4423 ( .A(n8641), .B(n8642), .C(n8643), .D(n8644), .Q(n8630) );
  NAND41 U4425 ( .A(n8669), .B(n8670), .C(n8671), .D(n8672), .Q(n8626) );
  NOR40 U4426 ( .A(n8673), .B(n8674), .C(n8675), .D(n8676), .Q(n8672) );
  NOR40 U4428 ( .A(n8677), .B(n8678), .C(n8679), .D(n8680), .Q(n8671) );
  NOR40 U4429 ( .A(n8681), .B(n8682), .C(n8683), .D(n8684), .Q(n8670) );
  NAND41 U4431 ( .A(n8713), .B(n8714), .C(n8715), .D(n8716), .Q(n8712) );
  NOR40 U4432 ( .A(n8717), .B(n8718), .C(n8719), .D(n8720), .Q(n8716) );
  NOR40 U4433 ( .A(n8721), .B(n8722), .C(n8723), .D(n8724), .Q(n8715) );
  NOR40 U4435 ( .A(n8725), .B(n8726), .C(n8727), .D(n8728), .Q(n8714) );
  NAND41 U4436 ( .A(n8753), .B(n8754), .C(n8755), .D(n8756), .Q(n8710) );
  NOR40 U4438 ( .A(n8757), .B(n8758), .C(n8759), .D(n8760), .Q(n8756) );
  NOR40 U4439 ( .A(n8761), .B(n8762), .C(n8763), .D(n8764), .Q(n8755) );
  NOR40 U4441 ( .A(n8765), .B(n8766), .C(n8767), .D(n8768), .Q(n8754) );
  NAND41 U4442 ( .A(n8799), .B(n8800), .C(n8801), .D(n8802), .Q(n8798) );
  NOR40 U4444 ( .A(n8803), .B(n8804), .C(n8805), .D(n8806), .Q(n8802) );
  NOR40 U4445 ( .A(n8807), .B(n8808), .C(n8809), .D(n8810), .Q(n8801) );
  NOR40 U4446 ( .A(n8811), .B(n8812), .C(n8813), .D(n8814), .Q(n8800) );
  NAND41 U4447 ( .A(n8839), .B(n8840), .C(n8841), .D(n8842), .Q(n8796) );
  NOR40 U4449 ( .A(n8843), .B(n8844), .C(n8845), .D(n8846), .Q(n8842) );
  NOR40 U4450 ( .A(n8847), .B(n8848), .C(n8849), .D(n8850), .Q(n8841) );
  NOR40 U4452 ( .A(n8851), .B(n8852), .C(n8853), .D(n8854), .Q(n8840) );
  NAND41 U4453 ( .A(n8883), .B(n8884), .C(n8885), .D(n8886), .Q(n8882) );
  NOR40 U4455 ( .A(n8887), .B(n8888), .C(n8889), .D(n8890), .Q(n8886) );
  NOR40 U4456 ( .A(n8891), .B(n8892), .C(n8893), .D(n8894), .Q(n8885) );
  NOR40 U4458 ( .A(n8895), .B(n8896), .C(n8897), .D(n8898), .Q(n8884) );
  NAND41 U4459 ( .A(n8923), .B(n8924), .C(n8925), .D(n8926), .Q(n8880) );
  NOR40 U4460 ( .A(n8927), .B(n8928), .C(n8929), .D(n8930), .Q(n8926) );
  NOR40 U4461 ( .A(n8931), .B(n8932), .C(n8933), .D(n8934), .Q(n8925) );
  NOR40 U4462 ( .A(n8935), .B(n8936), .C(n8937), .D(n8938), .Q(n8924) );
  NAND41 U4463 ( .A(n8969), .B(n8970), .C(n8971), .D(n8972), .Q(n8968) );
  NOR40 U4464 ( .A(n8973), .B(n8974), .C(n8975), .D(n8976), .Q(n8972) );
  NOR40 U4466 ( .A(n8977), .B(n8978), .C(n8979), .D(n8980), .Q(n8971) );
  NOR40 U4467 ( .A(n8981), .B(n8982), .C(n8983), .D(n8984), .Q(n8970) );
  NAND41 U4469 ( .A(n9009), .B(n9010), .C(n9011), .D(n9012), .Q(n8966) );
  NOR40 U4470 ( .A(n9013), .B(n9014), .C(n9015), .D(n9016), .Q(n9012) );
  NOR40 U4472 ( .A(n9017), .B(n9018), .C(n9019), .D(n9020), .Q(n9011) );
  NOR40 U4473 ( .A(n9021), .B(n9022), .C(n9023), .D(n9024), .Q(n9010) );
  NAND41 U4475 ( .A(n9053), .B(n9054), .C(n9055), .D(n9056), .Q(n9052) );
  NOR40 U4476 ( .A(n9057), .B(n9058), .C(n9059), .D(n9060), .Q(n9056) );
  NOR40 U4477 ( .A(n9061), .B(n9062), .C(n9063), .D(n9064), .Q(n9055) );
  NOR40 U4479 ( .A(n9065), .B(n9066), .C(n9067), .D(n9068), .Q(n9054) );
  NAND41 U4480 ( .A(n9093), .B(n9094), .C(n9095), .D(n9096), .Q(n9050) );
  NOR40 U4482 ( .A(n9097), .B(n9098), .C(n9099), .D(n9100), .Q(n9096) );
  NOR40 U4483 ( .A(n9101), .B(n9102), .C(n9103), .D(n9104), .Q(n9095) );
  NOR40 U4485 ( .A(n9105), .B(n9106), .C(n9107), .D(n9108), .Q(n9094) );
  NAND41 U4486 ( .A(n9139), .B(n9140), .C(n9141), .D(n9142), .Q(n9138) );
  NOR40 U4488 ( .A(n9143), .B(n9144), .C(n9145), .D(n9146), .Q(n9142) );
  NOR40 U4489 ( .A(n9147), .B(n9148), .C(n9149), .D(n9150), .Q(n9141) );
  NOR40 U4490 ( .A(n9151), .B(n9152), .C(n9153), .D(n9154), .Q(n9140) );
  NAND41 U4492 ( .A(n9179), .B(n9180), .C(n9181), .D(n9182), .Q(n9136) );
  NOR40 U4493 ( .A(n9183), .B(n9184), .C(n9185), .D(n9186), .Q(n9182) );
  NOR40 U4495 ( .A(n9187), .B(n9188), .C(n9189), .D(n9190), .Q(n9181) );
  NOR40 U4496 ( .A(n9191), .B(n9192), .C(n9193), .D(n9194), .Q(n9180) );
  NAND41 U4498 ( .A(n9223), .B(n9224), .C(n9225), .D(n9226), .Q(n9222) );
  NOR40 U4499 ( .A(n9227), .B(n9228), .C(n9229), .D(n9230), .Q(n9226) );
  NOR40 U4501 ( .A(n9231), .B(n9232), .C(n9233), .D(n9234), .Q(n9225) );
  NOR40 U4502 ( .A(n9235), .B(n9236), .C(n9237), .D(n9238), .Q(n9224) );
  NAND41 U4503 ( .A(n9263), .B(n9264), .C(n9265), .D(n9266), .Q(n9220) );
  NOR40 U4504 ( .A(n9267), .B(n9268), .C(n9269), .D(n9270), .Q(n9266) );
  NOR40 U4506 ( .A(n9271), .B(n9272), .C(n9273), .D(n9274), .Q(n9265) );
  NOR40 U4507 ( .A(n9275), .B(n9276), .C(n9277), .D(n9278), .Q(n9264) );
  NAND41 U4509 ( .A(n9309), .B(n9310), .C(n9311), .D(n9312), .Q(n9308) );
  NOR40 U4510 ( .A(n9313), .B(n9314), .C(n9315), .D(n9316), .Q(n9312) );
  NOR40 U4512 ( .A(n9317), .B(n9318), .C(n9319), .D(n9320), .Q(n9311) );
  NOR40 U4513 ( .A(n9321), .B(n9322), .C(n9323), .D(n9324), .Q(n9310) );
  NAND41 U4515 ( .A(n9349), .B(n9350), .C(n9351), .D(n9352), .Q(n9306) );
  NOR40 U4516 ( .A(n9353), .B(n9354), .C(n9355), .D(n9356), .Q(n9352) );
  NOR40 U4517 ( .A(n9357), .B(n9358), .C(n9359), .D(n9360), .Q(n9351) );
  NOR40 U4518 ( .A(n9361), .B(n9362), .C(n9363), .D(n9364), .Q(n9350) );
  NAND41 U4519 ( .A(n9393), .B(n9394), .C(n9395), .D(n9396), .Q(n9392) );
  NOR40 U4521 ( .A(n9397), .B(n9398), .C(n9399), .D(n9400), .Q(n9396) );
  NOR40 U4522 ( .A(n9401), .B(n9402), .C(n9403), .D(n9404), .Q(n9395) );
  NOR40 U4524 ( .A(n9405), .B(n9406), .C(n9407), .D(n9408), .Q(n9394) );
  NAND41 U4525 ( .A(n9433), .B(n9434), .C(n9435), .D(n9436), .Q(n9390) );
  NOR40 U4527 ( .A(n9437), .B(n9438), .C(n9439), .D(n9440), .Q(n9436) );
  NOR40 U4528 ( .A(n9441), .B(n9442), .C(n9443), .D(n9444), .Q(n9435) );
  NOR40 U4530 ( .A(n9445), .B(n9446), .C(n9447), .D(n9448), .Q(n9434) );
  NAND41 U4531 ( .A(n9479), .B(n9480), .C(n9481), .D(n9482), .Q(n9478) );
  NOR40 U4532 ( .A(n9483), .B(n9484), .C(n9485), .D(n9486), .Q(n9482) );
  NOR40 U4534 ( .A(n9487), .B(n9488), .C(n9489), .D(n9490), .Q(n9481) );
  NOR40 U4535 ( .A(n9491), .B(n9492), .C(n9493), .D(n9494), .Q(n9480) );
  NAND41 U4537 ( .A(n9519), .B(n9520), .C(n9521), .D(n9522), .Q(n9476) );
  NOR40 U4538 ( .A(n9523), .B(n9524), .C(n9525), .D(n9526), .Q(n9522) );
  NOR40 U4540 ( .A(n9527), .B(n9528), .C(n9529), .D(n9530), .Q(n9521) );
  NOR40 U4541 ( .A(n9531), .B(n9532), .C(n9533), .D(n9534), .Q(n9520) );
  NAND41 U4543 ( .A(n9563), .B(n9564), .C(n9565), .D(n9566), .Q(n9562) );
  NOR40 U4544 ( .A(n9567), .B(n9568), .C(n9569), .D(n9570), .Q(n9566) );
  NOR40 U4545 ( .A(n9571), .B(n9572), .C(n9573), .D(n9574), .Q(n9565) );
  NOR40 U4547 ( .A(n9575), .B(n9576), .C(n9577), .D(n9578), .Q(n9564) );
  NAND41 U4548 ( .A(n9603), .B(n9604), .C(n9605), .D(n9606), .Q(n9560) );
  NOR40 U4550 ( .A(n9607), .B(n9608), .C(n9609), .D(n9610), .Q(n9606) );
  NOR40 U4551 ( .A(n9611), .B(n9612), .C(n9613), .D(n9614), .Q(n9605) );
  NOR40 U4553 ( .A(n9615), .B(n9616), .C(n9617), .D(n9618), .Q(n9604) );
  NAND41 U4554 ( .A(n9649), .B(n9650), .C(n9651), .D(n9652), .Q(n9648) );
  NOR40 U4556 ( .A(n9653), .B(n9654), .C(n9655), .D(n9656), .Q(n9652) );
  NOR40 U4557 ( .A(n9657), .B(n9658), .C(n9659), .D(n9660), .Q(n9651) );
  NOR40 U4558 ( .A(n9661), .B(n9662), .C(n9663), .D(n9664), .Q(n9650) );
  NAND41 U4559 ( .A(n9689), .B(n9690), .C(n9691), .D(n9692), .Q(n9646) );
  NOR40 U4561 ( .A(n9693), .B(n9694), .C(n9695), .D(n9696), .Q(n9692) );
  NOR40 U4562 ( .A(n9697), .B(n9698), .C(n9699), .D(n9700), .Q(n9691) );
  NOR40 U4564 ( .A(n9701), .B(n9702), .C(n9703), .D(n9704), .Q(n9690) );
  NAND41 U4565 ( .A(n9733), .B(n9734), .C(n9735), .D(n9736), .Q(n9732) );
  NOR40 U4567 ( .A(n9737), .B(n9738), .C(n9739), .D(n9740), .Q(n9736) );
  NOR40 U4568 ( .A(n9741), .B(n9742), .C(n9743), .D(n9744), .Q(n9735) );
  NOR40 U4570 ( .A(n9745), .B(n9746), .C(n9747), .D(n9748), .Q(n9734) );
  NAND41 U4571 ( .A(n9773), .B(n9774), .C(n9775), .D(n9776), .Q(n9730) );
  NOR40 U4572 ( .A(n9777), .B(n9778), .C(n9779), .D(n9780), .Q(n9776) );
  NOR40 U4573 ( .A(n9781), .B(n9782), .C(n9783), .D(n9784), .Q(n9775) );
  NOR40 U4574 ( .A(n9785), .B(n9786), .C(n9787), .D(n9788), .Q(n9774) );
  NAND41 U4575 ( .A(n9819), .B(n9820), .C(n9821), .D(n9822), .Q(n9818) );
  NOR40 U4577 ( .A(n9823), .B(n9824), .C(n9825), .D(n9826), .Q(n9822) );
  NOR40 U4578 ( .A(n9827), .B(n9828), .C(n9829), .D(n9830), .Q(n9821) );
  NOR40 U4580 ( .A(n9831), .B(n9832), .C(n9833), .D(n9834), .Q(n9820) );
  NAND41 U4581 ( .A(n9859), .B(n9860), .C(n9861), .D(n9862), .Q(n9816) );
  NOR40 U4583 ( .A(n9863), .B(n9864), .C(n9865), .D(n9866), .Q(n9862) );
  NOR40 U4584 ( .A(n9867), .B(n9868), .C(n9869), .D(n9870), .Q(n9861) );
  NOR40 U4586 ( .A(n9871), .B(n9872), .C(n9873), .D(n9874), .Q(n9860) );
  NAND41 U4587 ( .A(n9903), .B(n9904), .C(n9905), .D(n9906), .Q(n9902) );
  NOR40 U4588 ( .A(n9907), .B(n9908), .C(n9909), .D(n9910), .Q(n9906) );
  NOR40 U4590 ( .A(n9911), .B(n9912), .C(n9913), .D(n9914), .Q(n9905) );
  NOR40 U4591 ( .A(n9915), .B(n9916), .C(n9917), .D(n9918), .Q(n9904) );
  NAND41 U4593 ( .A(n9943), .B(n9944), .C(n9945), .D(n9946), .Q(n9900) );
  NOR40 U4594 ( .A(n9947), .B(n9948), .C(n9949), .D(n9950), .Q(n9946) );
  NOR40 U4596 ( .A(n9951), .B(n9952), .C(n9953), .D(n9954), .Q(n9945) );
  NOR40 U4597 ( .A(n9955), .B(n9956), .C(n9957), .D(n9958), .Q(n9944) );
  NAND41 U4599 ( .A(n9989), .B(n9990), .C(n9991), .D(n9992), .Q(n9988) );
  NOR40 U4600 ( .A(n9993), .B(n9994), .C(n9995), .D(n9996), .Q(n9992) );
  NOR40 U4601 ( .A(n9997), .B(n9998), .C(n9999), .D(n10000), .Q(n9991) );
  NOR40 U4603 ( .A(n10001), .B(n10002), .C(n10003), .D(n10004), .Q(n9990) );
  NAND41 U4604 ( .A(n10029), .B(n10030), .C(n10031), .D(n10032), .Q(n9986) );
  NOR40 U4606 ( .A(n10033), .B(n10034), .C(n10035), .D(n10036), .Q(n10032) );
  NOR40 U4607 ( .A(n10037), .B(n10038), .C(n10039), .D(n10040), .Q(n10031) );
  NOR40 U4609 ( .A(n10041), .B(n10042), .C(n10043), .D(n10044), .Q(n10030) );
  NAND41 U4610 ( .A(n10073), .B(n10074), .C(n10075), .D(n10076), .Q(n10072) );
  NOR40 U4612 ( .A(n10077), .B(n10078), .C(n10079), .D(n10080), .Q(n10076) );
  NOR40 U4613 ( .A(n10081), .B(n10082), .C(n10083), .D(n10084), .Q(n10075) );
  NOR40 U4614 ( .A(n10085), .B(n10086), .C(n10087), .D(n10088), .Q(n10074) );
  NAND41 U4615 ( .A(n10113), .B(n10114), .C(n10115), .D(n10116), .Q(n10070) );
  NOR40 U4616 ( .A(n10117), .B(n10118), .C(n10119), .D(n10120), .Q(n10116) );
  NOR40 U4618 ( .A(n10121), .B(n10122), .C(n10123), .D(n10124), .Q(n10115) );
  NOR40 U4619 ( .A(n10125), .B(n10126), .C(n10127), .D(n10128), .Q(n10114) );
  NAND41 U4621 ( .A(n10159), .B(n10160), .C(n10161), .D(n10162), .Q(n10158) );
  NOR40 U4622 ( .A(n10163), .B(n10164), .C(n10165), .D(n10166), .Q(n10162) );
  NOR40 U4624 ( .A(n10167), .B(n10168), .C(n10169), .D(n10170), .Q(n10161) );
  NOR40 U4625 ( .A(n10171), .B(n10172), .C(n10173), .D(n10174), .Q(n10160) );
  NAND41 U4627 ( .A(n10199), .B(n10200), .C(n10201), .D(n10202), .Q(n10156) );
  NOR40 U4628 ( .A(n10203), .B(n10204), .C(n10205), .D(n10206), .Q(n10202) );
  NOR40 U4629 ( .A(n10207), .B(n10208), .C(n10209), .D(n10210), .Q(n10201) );
  NOR40 U4630 ( .A(n10211), .B(n10212), .C(n10213), .D(n10214), .Q(n10200) );
  NAND41 U4631 ( .A(n10243), .B(n10244), .C(n10245), .D(n10246), .Q(n10242) );
  NOR40 U4633 ( .A(n10247), .B(n10248), .C(n10249), .D(n10250), .Q(n10246) );
  NOR40 U4634 ( .A(n10251), .B(n10252), .C(n10253), .D(n10254), .Q(n10245) );
  NOR40 U4636 ( .A(n10255), .B(n10256), .C(n10257), .D(n10258), .Q(n10244) );
  NAND41 U4637 ( .A(n10283), .B(n10284), .C(n10285), .D(n10286), .Q(n10240) );
  NOR40 U4639 ( .A(n10287), .B(n10288), .C(n10289), .D(n10290), .Q(n10286) );
  NOR40 U4640 ( .A(n10291), .B(n10292), .C(n10293), .D(n10294), .Q(n10285) );
  NOR40 U4642 ( .A(n10295), .B(n10296), .C(n10297), .D(n10298), .Q(n10284) );
  NAND41 U4643 ( .A(n10329), .B(n10330), .C(n10331), .D(n10332), .Q(n10328) );
  NOR40 U4644 ( .A(n10333), .B(n10334), .C(n10335), .D(n10336), .Q(n10332) );
  NOR40 U4645 ( .A(n10337), .B(n10338), .C(n10339), .D(n10340), .Q(n10331) );
  NOR40 U4646 ( .A(n10341), .B(n10342), .C(n10343), .D(n10344), .Q(n10330) );
  NAND41 U4647 ( .A(n10369), .B(n10370), .C(n10371), .D(n10372), .Q(n10326) );
  NOR40 U4649 ( .A(n10373), .B(n10374), .C(n10375), .D(n10376), .Q(n10372) );
  NOR40 U4650 ( .A(n10377), .B(n10378), .C(n10379), .D(n10380), .Q(n10371) );
  NOR40 U4652 ( .A(n10381), .B(n10382), .C(n10383), .D(n10384), .Q(n10370) );
  NAND41 U4653 ( .A(n10413), .B(n10414), .C(n10415), .D(n10416), .Q(n10412) );
  NOR40 U4655 ( .A(n10417), .B(n10418), .C(n10419), .D(n10420), .Q(n10416) );
  NOR40 U4656 ( .A(n10421), .B(n10422), .C(n10423), .D(n10424), .Q(n10415) );
  NOR40 U4658 ( .A(n10425), .B(n10426), .C(n10427), .D(n10428), .Q(n10414) );
  NAND41 U4659 ( .A(n10453), .B(n10454), .C(n10455), .D(n10456), .Q(n10410) );
  NOR40 U4660 ( .A(n10457), .B(n10458), .C(n10459), .D(n10460), .Q(n10456) );
  NOR40 U4662 ( .A(n10461), .B(n10462), .C(n10463), .D(n10464), .Q(n10455) );
  NOR40 U4663 ( .A(n10465), .B(n10466), .C(n10467), .D(n10468), .Q(n10454) );
  NAND41 U4664 ( .A(n10499), .B(n10500), .C(n10501), .D(n10502), .Q(n10498) );
  NOR40 U4665 ( .A(n10503), .B(n10504), .C(n10505), .D(n10506), .Q(n10502) );
  NOR40 U4667 ( .A(n10507), .B(n10508), .C(n10509), .D(n10510), .Q(n10501) );
  NOR40 U4668 ( .A(n10511), .B(n10512), .C(n10513), .D(n10514), .Q(n10500) );
  NAND41 U4669 ( .A(n10539), .B(n10540), .C(n10541), .D(n10542), .Q(n10496) );
  NOR40 U4670 ( .A(n10543), .B(n10544), .C(n10545), .D(n10546), .Q(n10542) );
  NOR40 U4672 ( .A(n10547), .B(n10548), .C(n10549), .D(n10550), .Q(n10541) );
  NOR40 U4673 ( .A(n10551), .B(n10552), .C(n10553), .D(n10554), .Q(n10540) );
  NAND41 U4674 ( .A(n10583), .B(n10584), .C(n10585), .D(n10586), .Q(n10582) );
  NOR40 U4675 ( .A(n10587), .B(n10588), .C(n10589), .D(n10590), .Q(n10586) );
  NOR40 U4677 ( .A(n10591), .B(n10592), .C(n10593), .D(n10594), .Q(n10585) );
  NOR40 U4678 ( .A(n10595), .B(n10596), .C(n10597), .D(n10598), .Q(n10584) );
  NAND41 U4679 ( .A(n10623), .B(n10624), .C(n10625), .D(n10626), .Q(n10580) );
  NOR40 U4680 ( .A(n10627), .B(n10628), .C(n10629), .D(n10630), .Q(n10626) );
  NOR40 U4681 ( .A(n10631), .B(n10632), .C(n10633), .D(n10634), .Q(n10625) );
  NOR40 U4682 ( .A(n10635), .B(n10636), .C(n10637), .D(n10638), .Q(n10624) );
  NAND41 U4683 ( .A(n10669), .B(n10670), .C(n10671), .D(n10672), .Q(n10668) );
  NOR40 U4684 ( .A(n10673), .B(n10674), .C(n10675), .D(n10676), .Q(n10672) );
  NOR40 U4686 ( .A(n10677), .B(n10678), .C(n10679), .D(n10680), .Q(n10671) );
  NOR40 U4687 ( .A(n10681), .B(n10682), .C(n10683), .D(n10684), .Q(n10670) );
  NAND41 U4688 ( .A(n10716), .B(n10717), .C(n10718), .D(n10719), .Q(n10666) );
  NOR40 U4689 ( .A(n10720), .B(n10721), .C(n10722), .D(n10723), .Q(n10719) );
  NOR40 U4691 ( .A(n10724), .B(n10725), .C(n10726), .D(n10727), .Q(n10718) );
  NOR40 U4692 ( .A(n10728), .B(n10729), .C(n10730), .D(n10731), .Q(n10717) );
  NAND41 U4693 ( .A(n10766), .B(n10767), .C(n10768), .D(n10769), .Q(n10765) );
  NOR40 U4694 ( .A(n10770), .B(n10771), .C(n10772), .D(n10773), .Q(n10769) );
  NOR40 U4695 ( .A(n10774), .B(n10775), .C(n10776), .D(n10777), .Q(n10768) );
  NOR40 U4697 ( .A(n10778), .B(n10779), .C(n10780), .D(n10781), .Q(n10767) );
  NAND41 U4698 ( .A(n10811), .B(n10812), .C(n10813), .D(n10814), .Q(n10763) );
  NOR40 U4699 ( .A(n10815), .B(n10816), .C(n10817), .D(n10818), .Q(n10814) );
  NOR40 U4700 ( .A(n10819), .B(n10820), .C(n10821), .D(n10822), .Q(n10813) );
  NOR40 U4701 ( .A(n10823), .B(n10824), .C(n10825), .D(n10826), .Q(n10812) );
  NAND41 U4702 ( .A(n6659), .B(n6660), .C(n6661), .D(n6662), .Q(n6499) );
  NOR40 U4704 ( .A(n6663), .B(n6664), .C(n6665), .D(n6666), .Q(n6662) );
  NOR40 U4705 ( .A(n6675), .B(n6676), .C(n6677), .D(n6678), .Q(n6661) );
  NOR40 U4706 ( .A(n6687), .B(n6688), .C(n6689), .D(n6690), .Q(n6660) );
  NAND41 U4707 ( .A(n6989), .B(n6990), .C(n6991), .D(n6992), .Q(n6925) );
  NOR40 U4708 ( .A(n6993), .B(n6994), .C(n6995), .D(n6996), .Q(n6992) );
  NOR40 U4709 ( .A(n6997), .B(n6998), .C(n6999), .D(n7000), .Q(n6991) );
  NOR40 U4710 ( .A(n7001), .B(n7002), .C(n7003), .D(n7004), .Q(n6990) );
  NAND41 U4711 ( .A(n7159), .B(n7160), .C(n7161), .D(n7162), .Q(n7095) );
  NOR40 U4712 ( .A(n7163), .B(n7164), .C(n7165), .D(n7166), .Q(n7162) );
  NOR40 U4713 ( .A(n7167), .B(n7168), .C(n7169), .D(n7170), .Q(n7161) );
  NOR40 U4714 ( .A(n7171), .B(n7172), .C(n7173), .D(n7174), .Q(n7160) );
  NAND41 U4715 ( .A(n7329), .B(n7330), .C(n7331), .D(n7332), .Q(n7265) );
  NOR40 U4716 ( .A(n7333), .B(n7334), .C(n7335), .D(n7336), .Q(n7332) );
  NOR40 U4717 ( .A(n7337), .B(n7338), .C(n7339), .D(n7340), .Q(n7331) );
  NOR40 U4718 ( .A(n7341), .B(n7342), .C(n7343), .D(n7344), .Q(n7330) );
  NAND41 U4719 ( .A(n7499), .B(n7500), .C(n7501), .D(n7502), .Q(n7435) );
  NOR40 U4720 ( .A(n7503), .B(n7504), .C(n7505), .D(n7506), .Q(n7502) );
  NOR40 U4721 ( .A(n7507), .B(n7508), .C(n7509), .D(n7510), .Q(n7501) );
  NOR40 U4722 ( .A(n7511), .B(n7512), .C(n7513), .D(n7514), .Q(n7500) );
  NAND41 U4723 ( .A(n7669), .B(n7670), .C(n7671), .D(n7672), .Q(n7605) );
  NOR40 U4724 ( .A(n7673), .B(n7674), .C(n7675), .D(n7676), .Q(n7672) );
  NOR40 U4725 ( .A(n7677), .B(n7678), .C(n7679), .D(n7680), .Q(n7671) );
  NOR40 U4726 ( .A(n7681), .B(n7682), .C(n7683), .D(n7684), .Q(n7670) );
  NAND41 U4727 ( .A(n7839), .B(n7840), .C(n7841), .D(n7842), .Q(n7775) );
  NOR40 U4728 ( .A(n7843), .B(n7844), .C(n7845), .D(n7846), .Q(n7842) );
  NOR40 U4729 ( .A(n7847), .B(n7848), .C(n7849), .D(n7850), .Q(n7841) );
  NOR40 U4730 ( .A(n7851), .B(n7852), .C(n7853), .D(n7854), .Q(n7840) );
  NAND41 U4731 ( .A(n8009), .B(n8010), .C(n8011), .D(n8012), .Q(n7945) );
  NOR40 U4732 ( .A(n8013), .B(n8014), .C(n8015), .D(n8016), .Q(n8012) );
  NOR40 U4733 ( .A(n8017), .B(n8018), .C(n8019), .D(n8020), .Q(n8011) );
  NOR40 U4734 ( .A(n8021), .B(n8022), .C(n8023), .D(n8024), .Q(n8010) );
  NAND41 U4735 ( .A(n8179), .B(n8180), .C(n8181), .D(n8182), .Q(n8115) );
  NOR40 U4736 ( .A(n8183), .B(n8184), .C(n8185), .D(n8186), .Q(n8182) );
  NOR40 U4737 ( .A(n8187), .B(n8188), .C(n8189), .D(n8190), .Q(n8181) );
  NOR40 U4738 ( .A(n8191), .B(n8192), .C(n8193), .D(n8194), .Q(n8180) );
  NAND41 U4739 ( .A(n8349), .B(n8350), .C(n8351), .D(n8352), .Q(n8285) );
  NOR40 U4740 ( .A(n8353), .B(n8354), .C(n8355), .D(n8356), .Q(n8352) );
  NOR40 U4741 ( .A(n8357), .B(n8358), .C(n8359), .D(n8360), .Q(n8351) );
  NOR40 U4742 ( .A(n8361), .B(n8362), .C(n8363), .D(n8364), .Q(n8350) );
  NAND41 U4743 ( .A(n8519), .B(n8520), .C(n8521), .D(n8522), .Q(n8455) );
  NOR40 U4744 ( .A(n8523), .B(n8524), .C(n8525), .D(n8526), .Q(n8522) );
  NOR40 U4745 ( .A(n8527), .B(n8528), .C(n8529), .D(n8530), .Q(n8521) );
  NOR40 U4746 ( .A(n8531), .B(n8532), .C(n8533), .D(n8534), .Q(n8520) );
  NAND41 U4747 ( .A(n8689), .B(n8690), .C(n8691), .D(n8692), .Q(n8625) );
  NOR40 U4748 ( .A(n8693), .B(n8694), .C(n8695), .D(n8696), .Q(n8692) );
  NOR40 U4749 ( .A(n8697), .B(n8698), .C(n8699), .D(n8700), .Q(n8691) );
  NOR40 U4750 ( .A(n8701), .B(n8702), .C(n8703), .D(n8704), .Q(n8690) );
  NAND41 U4751 ( .A(n8859), .B(n8860), .C(n8861), .D(n8862), .Q(n8795) );
  NOR40 U4752 ( .A(n8863), .B(n8864), .C(n8865), .D(n8866), .Q(n8862) );
  NOR40 U4753 ( .A(n8867), .B(n8868), .C(n8869), .D(n8870), .Q(n8861) );
  NOR40 U4754 ( .A(n8871), .B(n8872), .C(n8873), .D(n8874), .Q(n8860) );
  NAND41 U4755 ( .A(n9029), .B(n9030), .C(n9031), .D(n9032), .Q(n8965) );
  NOR40 U4756 ( .A(n9033), .B(n9034), .C(n9035), .D(n9036), .Q(n9032) );
  NOR40 U4757 ( .A(n9037), .B(n9038), .C(n9039), .D(n9040), .Q(n9031) );
  NOR40 U4758 ( .A(n9041), .B(n9042), .C(n9043), .D(n9044), .Q(n9030) );
  NAND41 U4759 ( .A(n9199), .B(n9200), .C(n9201), .D(n9202), .Q(n9135) );
  NOR40 U4760 ( .A(n9203), .B(n9204), .C(n9205), .D(n9206), .Q(n9202) );
  NOR40 U4761 ( .A(n9207), .B(n9208), .C(n9209), .D(n9210), .Q(n9201) );
  NOR40 U4762 ( .A(n9211), .B(n9212), .C(n9213), .D(n9214), .Q(n9200) );
  NAND41 U4763 ( .A(n9369), .B(n9370), .C(n9371), .D(n9372), .Q(n9305) );
  NOR40 U4764 ( .A(n9373), .B(n9374), .C(n9375), .D(n9376), .Q(n9372) );
  NOR40 U4765 ( .A(n9377), .B(n9378), .C(n9379), .D(n9380), .Q(n9371) );
  NOR40 U4766 ( .A(n9381), .B(n9382), .C(n9383), .D(n9384), .Q(n9370) );
  NAND41 U4767 ( .A(n9539), .B(n9540), .C(n9541), .D(n9542), .Q(n9475) );
  NOR40 U4768 ( .A(n9543), .B(n9544), .C(n9545), .D(n9546), .Q(n9542) );
  NOR40 U4769 ( .A(n9547), .B(n9548), .C(n9549), .D(n9550), .Q(n9541) );
  NOR40 U4770 ( .A(n9551), .B(n9552), .C(n9553), .D(n9554), .Q(n9540) );
  NAND41 U4771 ( .A(n9709), .B(n9710), .C(n9711), .D(n9712), .Q(n9645) );
  NOR40 U4772 ( .A(n9713), .B(n9714), .C(n9715), .D(n9716), .Q(n9712) );
  NOR40 U4773 ( .A(n9717), .B(n9718), .C(n9719), .D(n9720), .Q(n9711) );
  NOR40 U4774 ( .A(n9721), .B(n9722), .C(n9723), .D(n9724), .Q(n9710) );
  NAND41 U4775 ( .A(n9879), .B(n9880), .C(n9881), .D(n9882), .Q(n9815) );
  NOR40 U4776 ( .A(n9883), .B(n9884), .C(n9885), .D(n9886), .Q(n9882) );
  NOR40 U4777 ( .A(n9887), .B(n9888), .C(n9889), .D(n9890), .Q(n9881) );
  NOR40 U4778 ( .A(n9891), .B(n9892), .C(n9893), .D(n9894), .Q(n9880) );
  NAND41 U4779 ( .A(n10049), .B(n10050), .C(n10051), .D(n10052), .Q(n9985) );
  NOR40 U4780 ( .A(n10053), .B(n10054), .C(n10055), .D(n10056), .Q(n10052) );
  NOR40 U4781 ( .A(n10057), .B(n10058), .C(n10059), .D(n10060), .Q(n10051) );
  NOR40 U4782 ( .A(n10061), .B(n10062), .C(n10063), .D(n10064), .Q(n10050) );
  NAND41 U4783 ( .A(n10219), .B(n10220), .C(n10221), .D(n10222), .Q(n10155) );
  NOR40 U4784 ( .A(n10223), .B(n10224), .C(n10225), .D(n10226), .Q(n10222) );
  NOR40 U4785 ( .A(n10227), .B(n10228), .C(n10229), .D(n10230), .Q(n10221) );
  NOR40 U4786 ( .A(n10231), .B(n10232), .C(n10233), .D(n10234), .Q(n10220) );
  NAND41 U4787 ( .A(n10389), .B(n10390), .C(n10391), .D(n10392), .Q(n10325) );
  NOR40 U4788 ( .A(n10393), .B(n10394), .C(n10395), .D(n10396), .Q(n10392) );
  NOR40 U4789 ( .A(n10397), .B(n10398), .C(n10399), .D(n10400), .Q(n10391) );
  NOR40 U4790 ( .A(n10401), .B(n10402), .C(n10403), .D(n10404), .Q(n10390) );
  NAND41 U4791 ( .A(n10559), .B(n10560), .C(n10561), .D(n10562), .Q(n10495) );
  NOR40 U4792 ( .A(n10563), .B(n10564), .C(n10565), .D(n10566), .Q(n10562) );
  NOR40 U4793 ( .A(n10567), .B(n10568), .C(n10569), .D(n10570), .Q(n10561) );
  NOR40 U4794 ( .A(n10571), .B(n10572), .C(n10573), .D(n10574), .Q(n10560) );
  NAND41 U4795 ( .A(n10740), .B(n10741), .C(n10742), .D(n10743), .Q(n10665) );
  NOR40 U4796 ( .A(n10744), .B(n10745), .C(n10746), .D(n10747), .Q(n10743) );
  NOR40 U4797 ( .A(n10748), .B(n10749), .C(n10750), .D(n10751), .Q(n10742) );
  NOR40 U4798 ( .A(n10752), .B(n10753), .C(n10754), .D(n10755), .Q(n10741) );
  NAND22 U4799 ( .A(n10864), .B(n10858), .Q(n10863) );
  NAND22 U4800 ( .A(n10709), .B(n10783), .Q(n10805) );
  NAND22 U4801 ( .A(n10715), .B(n10733), .Q(n10761) );
  NAND22 U4802 ( .A(n10715), .B(n10783), .Q(n10810) );
  NAND22 U4803 ( .A(n10687), .B(n10733), .Q(n10732) );
  NAND22 U4804 ( .A(n10687), .B(n10783), .Q(n10782) );
  NAND22 U4805 ( .A(n10733), .B(n10739), .Q(n10738) );
  NAND22 U4806 ( .A(n10828), .B(n10739), .Q(n10833) );
  NAND22 U4807 ( .A(n10686), .B(n10739), .Q(n10842) );
  NAND22 U4808 ( .A(n10686), .B(n10709), .Q(n10708) );
  NAND22 U4809 ( .A(n10686), .B(n10715), .Q(n10714) );
  NAND22 U4810 ( .A(n10686), .B(n10687), .Q(n10685) );
  NAND22 U4811 ( .A(n10828), .B(n10687), .Q(n10827) );
  NAND22 U4812 ( .A(n10828), .B(n10715), .Q(n10880) );
  NAND22 U4813 ( .A(n10828), .B(n10709), .Q(n10865) );
  NAND22 U4814 ( .A(n10853), .B(n10864), .Q(n10871) );
  NAND22 U4815 ( .A(n10853), .B(n10857), .Q(n10861) );
  NAND22 U4816 ( .A(n10857), .B(n10858), .Q(n10856) );
  NAND22 U4817 ( .A(n10874), .B(n10858), .Q(n10873) );
  NAND22 U4818 ( .A(n10852), .B(n10858), .Q(n10878) );
  NAND22 U4819 ( .A(n10852), .B(n10853), .Q(n10851) );
  NAND22 U4820 ( .A(n10874), .B(n10853), .Q(n10876) );
  NOR21 U4821 ( .A(n11343), .B(n11342), .Q(n10733) );
  NOR21 U4822 ( .A(n11323), .B(n11322), .Q(n10857) );
  NAND22 U4823 ( .A(n6497), .B(n6498), .Q(N814) );
  NOR40 U4824 ( .A(n6711), .B(n6712), .C(n6713), .D(n6714), .Q(n6497) );
  NOR40 U4825 ( .A(n6499), .B(n6500), .C(n6501), .D(n6502), .Q(n6498) );
  NAND41 U4826 ( .A(n6871), .B(n6872), .C(n6873), .D(n6874), .Q(n6711) );
  NAND22 U4827 ( .A(n6923), .B(n6924), .Q(N813) );
  NOR40 U4828 ( .A(n7009), .B(n7010), .C(n7011), .D(n7012), .Q(n6923) );
  NOR40 U4829 ( .A(n6925), .B(n6926), .C(n6927), .D(n6928), .Q(n6924) );
  NAND41 U4830 ( .A(n7073), .B(n7074), .C(n7075), .D(n7076), .Q(n7009) );
  NAND22 U4831 ( .A(n7093), .B(n7094), .Q(N812) );
  NOR40 U4832 ( .A(n7179), .B(n7180), .C(n7181), .D(n7182), .Q(n7093) );
  NOR40 U4833 ( .A(n7095), .B(n7096), .C(n7097), .D(n7098), .Q(n7094) );
  NAND41 U4834 ( .A(n7243), .B(n7244), .C(n7245), .D(n7246), .Q(n7179) );
  NAND22 U4835 ( .A(n7263), .B(n7264), .Q(N811) );
  NOR40 U4836 ( .A(n7349), .B(n7350), .C(n7351), .D(n7352), .Q(n7263) );
  NOR40 U4837 ( .A(n7265), .B(n7266), .C(n7267), .D(n7268), .Q(n7264) );
  NAND41 U4838 ( .A(n7413), .B(n7414), .C(n7415), .D(n7416), .Q(n7349) );
  NAND22 U4839 ( .A(n7433), .B(n7434), .Q(N810) );
  NOR40 U4840 ( .A(n7519), .B(n7520), .C(n7521), .D(n7522), .Q(n7433) );
  NOR40 U4841 ( .A(n7435), .B(n7436), .C(n7437), .D(n7438), .Q(n7434) );
  NAND41 U4842 ( .A(n7583), .B(n7584), .C(n7585), .D(n7586), .Q(n7519) );
  NAND22 U4843 ( .A(n7603), .B(n7604), .Q(N809) );
  NOR40 U4844 ( .A(n7689), .B(n7690), .C(n7691), .D(n7692), .Q(n7603) );
  NOR40 U4845 ( .A(n7605), .B(n7606), .C(n7607), .D(n7608), .Q(n7604) );
  NAND41 U4846 ( .A(n7753), .B(n7754), .C(n7755), .D(n7756), .Q(n7689) );
  NAND22 U4847 ( .A(n7773), .B(n7774), .Q(N808) );
  NOR40 U4848 ( .A(n7859), .B(n7860), .C(n7861), .D(n7862), .Q(n7773) );
  NOR40 U4849 ( .A(n7775), .B(n7776), .C(n7777), .D(n7778), .Q(n7774) );
  NAND41 U4850 ( .A(n7923), .B(n7924), .C(n7925), .D(n7926), .Q(n7859) );
  NAND22 U4851 ( .A(n7943), .B(n7944), .Q(N807) );
  NOR40 U4852 ( .A(n8029), .B(n8030), .C(n8031), .D(n8032), .Q(n7943) );
  NOR40 U4853 ( .A(n7945), .B(n7946), .C(n7947), .D(n7948), .Q(n7944) );
  NAND41 U4854 ( .A(n8093), .B(n8094), .C(n8095), .D(n8096), .Q(n8029) );
  NAND22 U4855 ( .A(n8113), .B(n8114), .Q(N806) );
  NOR40 U4856 ( .A(n8199), .B(n8200), .C(n8201), .D(n8202), .Q(n8113) );
  NOR40 U4857 ( .A(n8115), .B(n8116), .C(n8117), .D(n8118), .Q(n8114) );
  NAND41 U4858 ( .A(n8263), .B(n8264), .C(n8265), .D(n8266), .Q(n8199) );
  NAND22 U4859 ( .A(n8283), .B(n8284), .Q(N805) );
  NOR40 U4860 ( .A(n8369), .B(n8370), .C(n8371), .D(n8372), .Q(n8283) );
  NOR40 U4861 ( .A(n8285), .B(n8286), .C(n8287), .D(n8288), .Q(n8284) );
  NAND41 U4862 ( .A(n8433), .B(n8434), .C(n8435), .D(n8436), .Q(n8369) );
  NAND22 U4863 ( .A(n8453), .B(n8454), .Q(N804) );
  NOR40 U4864 ( .A(n8539), .B(n8540), .C(n8541), .D(n8542), .Q(n8453) );
  NOR40 U4865 ( .A(n8455), .B(n8456), .C(n8457), .D(n8458), .Q(n8454) );
  NAND41 U4866 ( .A(n8603), .B(n8604), .C(n8605), .D(n8606), .Q(n8539) );
  NAND22 U4867 ( .A(n8623), .B(n8624), .Q(N803) );
  NOR40 U4868 ( .A(n8709), .B(n8710), .C(n8711), .D(n8712), .Q(n8623) );
  NOR40 U4869 ( .A(n8625), .B(n8626), .C(n8627), .D(n8628), .Q(n8624) );
  NAND41 U4870 ( .A(n8773), .B(n8774), .C(n8775), .D(n8776), .Q(n8709) );
  NAND22 U4871 ( .A(n8793), .B(n8794), .Q(N802) );
  NOR40 U4872 ( .A(n8879), .B(n8880), .C(n8881), .D(n8882), .Q(n8793) );
  NOR40 U4873 ( .A(n8795), .B(n8796), .C(n8797), .D(n8798), .Q(n8794) );
  NAND41 U4874 ( .A(n8943), .B(n8944), .C(n8945), .D(n8946), .Q(n8879) );
  NAND22 U4875 ( .A(n8963), .B(n8964), .Q(N801) );
  NOR40 U4876 ( .A(n9049), .B(n9050), .C(n9051), .D(n9052), .Q(n8963) );
  NOR40 U4877 ( .A(n8965), .B(n8966), .C(n8967), .D(n8968), .Q(n8964) );
  NAND41 U4878 ( .A(n9113), .B(n9114), .C(n9115), .D(n9116), .Q(n9049) );
  NAND22 U4879 ( .A(n9133), .B(n9134), .Q(N800) );
  NOR40 U4880 ( .A(n9219), .B(n9220), .C(n9221), .D(n9222), .Q(n9133) );
  NOR40 U4881 ( .A(n9135), .B(n9136), .C(n9137), .D(n9138), .Q(n9134) );
  NAND41 U4882 ( .A(n9283), .B(n9284), .C(n9285), .D(n9286), .Q(n9219) );
  NAND22 U4883 ( .A(n9303), .B(n9304), .Q(N799) );
  NOR40 U4884 ( .A(n9389), .B(n9390), .C(n9391), .D(n9392), .Q(n9303) );
  NOR40 U4885 ( .A(n9305), .B(n9306), .C(n9307), .D(n9308), .Q(n9304) );
  NAND41 U4886 ( .A(n9453), .B(n9454), .C(n9455), .D(n9456), .Q(n9389) );
  NAND22 U4887 ( .A(n9473), .B(n9474), .Q(N798) );
  NOR40 U4888 ( .A(n9559), .B(n9560), .C(n9561), .D(n9562), .Q(n9473) );
  NOR40 U4889 ( .A(n9475), .B(n9476), .C(n9477), .D(n9478), .Q(n9474) );
  NAND41 U4890 ( .A(n9623), .B(n9624), .C(n9625), .D(n9626), .Q(n9559) );
  NAND22 U4891 ( .A(n9643), .B(n9644), .Q(N797) );
  NOR40 U4892 ( .A(n9729), .B(n9730), .C(n9731), .D(n9732), .Q(n9643) );
  NOR40 U4893 ( .A(n9645), .B(n9646), .C(n9647), .D(n9648), .Q(n9644) );
  NAND41 U4894 ( .A(n9793), .B(n9794), .C(n9795), .D(n9796), .Q(n9729) );
  NAND22 U4895 ( .A(n9813), .B(n9814), .Q(N796) );
  NOR40 U4896 ( .A(n9899), .B(n9900), .C(n9901), .D(n9902), .Q(n9813) );
  NOR40 U4897 ( .A(n9815), .B(n9816), .C(n9817), .D(n9818), .Q(n9814) );
  NAND41 U4898 ( .A(n9963), .B(n9964), .C(n9965), .D(n9966), .Q(n9899) );
  NAND22 U4899 ( .A(n9983), .B(n9984), .Q(N795) );
  NOR40 U4900 ( .A(n10069), .B(n10070), .C(n10071), .D(n10072), .Q(n9983) );
  NOR40 U4901 ( .A(n9985), .B(n9986), .C(n9987), .D(n9988), .Q(n9984) );
  NAND41 U4902 ( .A(n10133), .B(n10134), .C(n10135), .D(n10136), .Q(n10069) );
  NAND22 U4903 ( .A(n10153), .B(n10154), .Q(N794) );
  NOR40 U4904 ( .A(n10239), .B(n10240), .C(n10241), .D(n10242), .Q(n10153) );
  NOR40 U4905 ( .A(n10155), .B(n10156), .C(n10157), .D(n10158), .Q(n10154) );
  NAND41 U4906 ( .A(n10303), .B(n10304), .C(n10305), .D(n10306), .Q(n10239) );
  NAND22 U4907 ( .A(n10323), .B(n10324), .Q(N793) );
  NOR40 U4908 ( .A(n10409), .B(n10410), .C(n10411), .D(n10412), .Q(n10323) );
  NOR40 U4909 ( .A(n10325), .B(n10326), .C(n10327), .D(n10328), .Q(n10324) );
  NAND41 U4910 ( .A(n10473), .B(n10474), .C(n10475), .D(n10476), .Q(n10409) );
  NAND22 U4911 ( .A(n10493), .B(n10494), .Q(N792) );
  NOR40 U4912 ( .A(n10579), .B(n10580), .C(n10581), .D(n10582), .Q(n10493) );
  NOR40 U4913 ( .A(n10495), .B(n10496), .C(n10497), .D(n10498), .Q(n10494) );
  NAND41 U4914 ( .A(n10643), .B(n10644), .C(n10645), .D(n10646), .Q(n10579) );
  NAND22 U4915 ( .A(n10663), .B(n10664), .Q(N791) );
  NOR40 U4916 ( .A(n10762), .B(n10763), .C(n10764), .D(n10765), .Q(n10663) );
  NOR40 U4917 ( .A(n10665), .B(n10666), .C(n10667), .D(n10668), .Q(n10664) );
  NAND41 U4918 ( .A(n10834), .B(n10835), .C(n10836), .D(n10837), .Q(n10762) );
  NOR21 U4919 ( .A(n11351), .B(waddr_6), .Q(n6312) );
  NOR21 U4920 ( .A(n11348), .B(waddr_5), .Q(n6255) );
  NOR21 U4921 ( .A(n11349), .B(waddr_4), .Q(n6274) );
  NOR21 U4922 ( .A(n11350), .B(waddr_7), .Q(n6235) );
  NOR21 U4923 ( .A(waddr_7), .B(waddr_6), .Q(n6438) );
  INV3 U4924 ( .A(waddr_1), .Q(n11345) );
  INV3 U4925 ( .A(waddr_0), .Q(n11344) );
  NAND31 U4926 ( .A(wreq), .B(n6438), .C(n6234), .Q(n6420) );
  NAND31 U4927 ( .A(n6381), .B(wreq), .C(n6234), .Q(n6365) );
  NAND31 U4928 ( .A(n6234), .B(wreq), .C(n6312), .Q(n6296) );
  NAND31 U4929 ( .A(n6255), .B(wreq), .C(n6312), .Q(n6314) );
  NAND31 U4930 ( .A(n6274), .B(wreq), .C(n6312), .Q(n6331) );
  NAND31 U4931 ( .A(wreq), .B(n6294), .C(n6312), .Q(n6348) );
  NAND31 U4932 ( .A(wreq), .B(n6438), .C(n6255), .Q(n6440) );
  NAND31 U4933 ( .A(n6235), .B(wreq), .C(n6255), .Q(n6237) );
  NAND31 U4934 ( .A(n6381), .B(wreq), .C(n6255), .Q(n6383) );
  NAND31 U4935 ( .A(wreq), .B(n6438), .C(n6274), .Q(n6458) );
  NAND31 U4936 ( .A(n6235), .B(wreq), .C(n6274), .Q(n6257) );
  NAND31 U4937 ( .A(n6381), .B(wreq), .C(n6274), .Q(n6400) );
  NAND31 U4938 ( .A(n6234), .B(wreq), .C(n6235), .Q(n6202) );
  NAND31 U4939 ( .A(wreq), .B(n6294), .C(n6235), .Q(n6276) );
  INV3 U4940 ( .A(waddr_5), .Q(n11349) );
  INV3 U4941 ( .A(waddr_3), .Q(n11347) );
  NAND31 U4942 ( .A(wreq), .B(n6294), .C(n6381), .Q(n6222) );
  INV3 U4943 ( .A(waddr_7), .Q(n11351) );
  INV3 U4944 ( .A(waddr_6), .Q(n11350) );
  INV3 U4945 ( .A(waddr_4), .Q(n11348) );
  INV3 U4946 ( .A(waddr_2), .Q(n11346) );
  NAND31 U4947 ( .A(n6294), .B(n6438), .C(wreq), .Q(n6197) );
  NOR21 U4948 ( .A(n11321), .B(raddr_0), .Q(n10853) );
  NOR21 U4949 ( .A(n11312), .B(raddr_1), .Q(n10855) );
  NOR21 U4950 ( .A(n11341), .B(raddr_4), .Q(n10715) );
  NOR21 U4951 ( .A(n11332), .B(raddr_5), .Q(n10687) );
  NOR40 U4952 ( .A(n6595), .B(n6596), .C(n6597), .D(n6598), .Q(n6555) );
  NOR40 U4953 ( .A(n6543), .B(n6544), .C(n6545), .D(n6546), .Q(n6503) );
  NOR40 U4954 ( .A(n6647), .B(n6648), .C(n6649), .D(n6650), .Q(n6607) );
  NOR40 U4955 ( .A(n6699), .B(n6700), .C(n6701), .D(n6702), .Q(n6659) );
  NOR40 U4956 ( .A(n6807), .B(n6808), .C(n6809), .D(n6810), .Q(n6767) );
  NOR40 U4957 ( .A(n6755), .B(n6756), .C(n6757), .D(n6758), .Q(n6715) );
  NOR40 U4958 ( .A(n6859), .B(n6860), .C(n6861), .D(n6862), .Q(n6819) );
  NOR40 U4959 ( .A(n6911), .B(n6912), .C(n6913), .D(n6914), .Q(n6871) );
  NOR40 U4960 ( .A(n6965), .B(n6966), .C(n6967), .D(n6968), .Q(n6949) );
  NOR40 U4961 ( .A(n6945), .B(n6946), .C(n6947), .D(n6948), .Q(n6929) );
  NOR40 U4962 ( .A(n6985), .B(n6986), .C(n6987), .D(n6988), .Q(n6969) );
  NOR40 U4963 ( .A(n7005), .B(n7006), .C(n7007), .D(n7008), .Q(n6989) );
  NOR40 U4964 ( .A(n7049), .B(n7050), .C(n7051), .D(n7052), .Q(n7033) );
  NOR40 U4965 ( .A(n7029), .B(n7030), .C(n7031), .D(n7032), .Q(n7013) );
  NOR40 U4966 ( .A(n7069), .B(n7070), .C(n7071), .D(n7072), .Q(n7053) );
  NOR40 U4967 ( .A(n7089), .B(n7090), .C(n7091), .D(n7092), .Q(n7073) );
  NOR40 U4968 ( .A(n7135), .B(n7136), .C(n7137), .D(n7138), .Q(n7119) );
  NOR40 U4969 ( .A(n7115), .B(n7116), .C(n7117), .D(n7118), .Q(n7099) );
  NOR40 U4970 ( .A(n7155), .B(n7156), .C(n7157), .D(n7158), .Q(n7139) );
  NOR40 U4971 ( .A(n7175), .B(n7176), .C(n7177), .D(n7178), .Q(n7159) );
  NOR40 U4972 ( .A(n7219), .B(n7220), .C(n7221), .D(n7222), .Q(n7203) );
  NOR40 U4973 ( .A(n7199), .B(n7200), .C(n7201), .D(n7202), .Q(n7183) );
  NOR40 U4974 ( .A(n7239), .B(n7240), .C(n7241), .D(n7242), .Q(n7223) );
  NOR40 U4975 ( .A(n7259), .B(n7260), .C(n7261), .D(n7262), .Q(n7243) );
  NOR40 U4976 ( .A(n7305), .B(n7306), .C(n7307), .D(n7308), .Q(n7289) );
  NOR40 U4977 ( .A(n7285), .B(n7286), .C(n7287), .D(n7288), .Q(n7269) );
  NOR40 U4978 ( .A(n7325), .B(n7326), .C(n7327), .D(n7328), .Q(n7309) );
  NOR40 U4979 ( .A(n7345), .B(n7346), .C(n7347), .D(n7348), .Q(n7329) );
  NOR40 U4980 ( .A(n7389), .B(n7390), .C(n7391), .D(n7392), .Q(n7373) );
  NOR40 U4981 ( .A(n7369), .B(n7370), .C(n7371), .D(n7372), .Q(n7353) );
  NOR40 U4982 ( .A(n7409), .B(n7410), .C(n7411), .D(n7412), .Q(n7393) );
  NOR40 U4983 ( .A(n7429), .B(n7430), .C(n7431), .D(n7432), .Q(n7413) );
  NOR40 U4984 ( .A(n7475), .B(n7476), .C(n7477), .D(n7478), .Q(n7459) );
  NOR40 U4985 ( .A(n7455), .B(n7456), .C(n7457), .D(n7458), .Q(n7439) );
  NOR40 U4986 ( .A(n7495), .B(n7496), .C(n7497), .D(n7498), .Q(n7479) );
  NOR40 U4987 ( .A(n7515), .B(n7516), .C(n7517), .D(n7518), .Q(n7499) );
  NOR40 U4988 ( .A(n7559), .B(n7560), .C(n7561), .D(n7562), .Q(n7543) );
  NOR40 U4989 ( .A(n7539), .B(n7540), .C(n7541), .D(n7542), .Q(n7523) );
  NOR40 U4990 ( .A(n7579), .B(n7580), .C(n7581), .D(n7582), .Q(n7563) );
  NOR40 U4991 ( .A(n7599), .B(n7600), .C(n7601), .D(n7602), .Q(n7583) );
  NOR40 U4992 ( .A(n7645), .B(n7646), .C(n7647), .D(n7648), .Q(n7629) );
  NOR40 U4993 ( .A(n7625), .B(n7626), .C(n7627), .D(n7628), .Q(n7609) );
  NOR40 U4994 ( .A(n7665), .B(n7666), .C(n7667), .D(n7668), .Q(n7649) );
  NOR40 U4995 ( .A(n7685), .B(n7686), .C(n7687), .D(n7688), .Q(n7669) );
  NOR40 U4996 ( .A(n7729), .B(n7730), .C(n7731), .D(n7732), .Q(n7713) );
  NOR40 U4997 ( .A(n7709), .B(n7710), .C(n7711), .D(n7712), .Q(n7693) );
  NOR40 U4998 ( .A(n7749), .B(n7750), .C(n7751), .D(n7752), .Q(n7733) );
  NOR40 U4999 ( .A(n7769), .B(n7770), .C(n7771), .D(n7772), .Q(n7753) );
  NOR40 U5000 ( .A(n7815), .B(n7816), .C(n7817), .D(n7818), .Q(n7799) );
  NOR40 U5001 ( .A(n7795), .B(n7796), .C(n7797), .D(n7798), .Q(n7779) );
  NOR40 U5002 ( .A(n7835), .B(n7836), .C(n7837), .D(n7838), .Q(n7819) );
  NOR40 U5003 ( .A(n7855), .B(n7856), .C(n7857), .D(n7858), .Q(n7839) );
  NOR40 U5004 ( .A(n7899), .B(n7900), .C(n7901), .D(n7902), .Q(n7883) );
  NOR40 U5005 ( .A(n7879), .B(n7880), .C(n7881), .D(n7882), .Q(n7863) );
  NOR40 U5006 ( .A(n7919), .B(n7920), .C(n7921), .D(n7922), .Q(n7903) );
  NOR40 U5007 ( .A(n7939), .B(n7940), .C(n7941), .D(n7942), .Q(n7923) );
  NOR40 U5008 ( .A(n7985), .B(n7986), .C(n7987), .D(n7988), .Q(n7969) );
  NOR40 U5009 ( .A(n7965), .B(n7966), .C(n7967), .D(n7968), .Q(n7949) );
  NOR40 U5010 ( .A(n8005), .B(n8006), .C(n8007), .D(n8008), .Q(n7989) );
  NOR40 U5011 ( .A(n8025), .B(n8026), .C(n8027), .D(n8028), .Q(n8009) );
  NOR40 U5012 ( .A(n8069), .B(n8070), .C(n8071), .D(n8072), .Q(n8053) );
  NOR40 U5013 ( .A(n8049), .B(n8050), .C(n8051), .D(n8052), .Q(n8033) );
  NOR40 U5014 ( .A(n8089), .B(n8090), .C(n8091), .D(n8092), .Q(n8073) );
  NOR40 U5015 ( .A(n8109), .B(n8110), .C(n8111), .D(n8112), .Q(n8093) );
  NOR40 U5016 ( .A(n8155), .B(n8156), .C(n8157), .D(n8158), .Q(n8139) );
  NOR40 U5017 ( .A(n8135), .B(n8136), .C(n8137), .D(n8138), .Q(n8119) );
  NOR40 U5018 ( .A(n8175), .B(n8176), .C(n8177), .D(n8178), .Q(n8159) );
  NOR40 U5019 ( .A(n8195), .B(n8196), .C(n8197), .D(n8198), .Q(n8179) );
  NOR40 U5020 ( .A(n8239), .B(n8240), .C(n8241), .D(n8242), .Q(n8223) );
  NOR40 U5021 ( .A(n8219), .B(n8220), .C(n8221), .D(n8222), .Q(n8203) );
  NOR40 U5022 ( .A(n8259), .B(n8260), .C(n8261), .D(n8262), .Q(n8243) );
  NOR40 U5023 ( .A(n8279), .B(n8280), .C(n8281), .D(n8282), .Q(n8263) );
  NOR40 U5024 ( .A(n8325), .B(n8326), .C(n8327), .D(n8328), .Q(n8309) );
  NOR40 U5025 ( .A(n8305), .B(n8306), .C(n8307), .D(n8308), .Q(n8289) );
  NOR40 U5026 ( .A(n8345), .B(n8346), .C(n8347), .D(n8348), .Q(n8329) );
  NOR40 U5027 ( .A(n8365), .B(n8366), .C(n8367), .D(n8368), .Q(n8349) );
  NOR40 U5028 ( .A(n8409), .B(n8410), .C(n8411), .D(n8412), .Q(n8393) );
  NOR40 U5029 ( .A(n8389), .B(n8390), .C(n8391), .D(n8392), .Q(n8373) );
  NOR40 U5030 ( .A(n8429), .B(n8430), .C(n8431), .D(n8432), .Q(n8413) );
  NOR40 U5031 ( .A(n8449), .B(n8450), .C(n8451), .D(n8452), .Q(n8433) );
  NOR40 U5032 ( .A(n8495), .B(n8496), .C(n8497), .D(n8498), .Q(n8479) );
  NOR40 U5033 ( .A(n8475), .B(n8476), .C(n8477), .D(n8478), .Q(n8459) );
  NOR40 U5034 ( .A(n8515), .B(n8516), .C(n8517), .D(n8518), .Q(n8499) );
  NOR40 U5035 ( .A(n8535), .B(n8536), .C(n8537), .D(n8538), .Q(n8519) );
  NOR40 U5036 ( .A(n8579), .B(n8580), .C(n8581), .D(n8582), .Q(n8563) );
  NOR40 U5037 ( .A(n8559), .B(n8560), .C(n8561), .D(n8562), .Q(n8543) );
  NOR40 U5038 ( .A(n8599), .B(n8600), .C(n8601), .D(n8602), .Q(n8583) );
  NOR40 U5039 ( .A(n8619), .B(n8620), .C(n8621), .D(n8622), .Q(n8603) );
  NOR40 U5040 ( .A(n8665), .B(n8666), .C(n8667), .D(n8668), .Q(n8649) );
  NOR40 U5041 ( .A(n8645), .B(n8646), .C(n8647), .D(n8648), .Q(n8629) );
  NOR40 U5042 ( .A(n8685), .B(n8686), .C(n8687), .D(n8688), .Q(n8669) );
  NOR40 U5043 ( .A(n8705), .B(n8706), .C(n8707), .D(n8708), .Q(n8689) );
  NOR40 U5044 ( .A(n8749), .B(n8750), .C(n8751), .D(n8752), .Q(n8733) );
  NOR40 U5045 ( .A(n8729), .B(n8730), .C(n8731), .D(n8732), .Q(n8713) );
  NOR40 U5046 ( .A(n8769), .B(n8770), .C(n8771), .D(n8772), .Q(n8753) );
  NOR40 U5047 ( .A(n8789), .B(n8790), .C(n8791), .D(n8792), .Q(n8773) );
  NOR40 U5048 ( .A(n8835), .B(n8836), .C(n8837), .D(n8838), .Q(n8819) );
  NOR40 U5049 ( .A(n8815), .B(n8816), .C(n8817), .D(n8818), .Q(n8799) );
  NOR40 U5050 ( .A(n8855), .B(n8856), .C(n8857), .D(n8858), .Q(n8839) );
  NOR40 U5051 ( .A(n8875), .B(n8876), .C(n8877), .D(n8878), .Q(n8859) );
  NOR40 U5052 ( .A(n8919), .B(n8920), .C(n8921), .D(n8922), .Q(n8903) );
  NOR40 U5053 ( .A(n8899), .B(n8900), .C(n8901), .D(n8902), .Q(n8883) );
  NOR40 U5054 ( .A(n8939), .B(n8940), .C(n8941), .D(n8942), .Q(n8923) );
  NOR40 U5055 ( .A(n8959), .B(n8960), .C(n8961), .D(n8962), .Q(n8943) );
  NOR40 U5056 ( .A(n9005), .B(n9006), .C(n9007), .D(n9008), .Q(n8989) );
  NOR40 U5057 ( .A(n8985), .B(n8986), .C(n8987), .D(n8988), .Q(n8969) );
  NOR40 U5058 ( .A(n9025), .B(n9026), .C(n9027), .D(n9028), .Q(n9009) );
  NOR40 U5059 ( .A(n9045), .B(n9046), .C(n9047), .D(n9048), .Q(n9029) );
  NOR40 U5060 ( .A(n9089), .B(n9090), .C(n9091), .D(n9092), .Q(n9073) );
  NOR40 U5061 ( .A(n9069), .B(n9070), .C(n9071), .D(n9072), .Q(n9053) );
  NOR40 U5062 ( .A(n9109), .B(n9110), .C(n9111), .D(n9112), .Q(n9093) );
  NOR40 U5063 ( .A(n9129), .B(n9130), .C(n9131), .D(n9132), .Q(n9113) );
  NOR40 U5064 ( .A(n9175), .B(n9176), .C(n9177), .D(n9178), .Q(n9159) );
  NOR40 U5065 ( .A(n9155), .B(n9156), .C(n9157), .D(n9158), .Q(n9139) );
  NOR40 U5066 ( .A(n9195), .B(n9196), .C(n9197), .D(n9198), .Q(n9179) );
  NOR40 U5067 ( .A(n9215), .B(n9216), .C(n9217), .D(n9218), .Q(n9199) );
  NOR40 U5068 ( .A(n9259), .B(n9260), .C(n9261), .D(n9262), .Q(n9243) );
  NOR40 U5069 ( .A(n9239), .B(n9240), .C(n9241), .D(n9242), .Q(n9223) );
  NOR40 U5070 ( .A(n9279), .B(n9280), .C(n9281), .D(n9282), .Q(n9263) );
  NOR40 U5071 ( .A(n9299), .B(n9300), .C(n9301), .D(n9302), .Q(n9283) );
  NOR40 U5072 ( .A(n9345), .B(n9346), .C(n9347), .D(n9348), .Q(n9329) );
  NOR40 U5073 ( .A(n9325), .B(n9326), .C(n9327), .D(n9328), .Q(n9309) );
  NOR40 U5074 ( .A(n9365), .B(n9366), .C(n9367), .D(n9368), .Q(n9349) );
  NOR40 U5075 ( .A(n9385), .B(n9386), .C(n9387), .D(n9388), .Q(n9369) );
  NOR40 U5076 ( .A(n9429), .B(n9430), .C(n9431), .D(n9432), .Q(n9413) );
  NOR40 U5077 ( .A(n9409), .B(n9410), .C(n9411), .D(n9412), .Q(n9393) );
  NOR40 U5078 ( .A(n9449), .B(n9450), .C(n9451), .D(n9452), .Q(n9433) );
  NOR40 U5079 ( .A(n9469), .B(n9470), .C(n9471), .D(n9472), .Q(n9453) );
  NOR40 U5080 ( .A(n9515), .B(n9516), .C(n9517), .D(n9518), .Q(n9499) );
  NOR40 U5081 ( .A(n9495), .B(n9496), .C(n9497), .D(n9498), .Q(n9479) );
  NOR40 U5082 ( .A(n9535), .B(n9536), .C(n9537), .D(n9538), .Q(n9519) );
  NOR40 U5083 ( .A(n9555), .B(n9556), .C(n9557), .D(n9558), .Q(n9539) );
  NOR40 U5084 ( .A(n9599), .B(n9600), .C(n9601), .D(n9602), .Q(n9583) );
  NOR40 U5085 ( .A(n9579), .B(n9580), .C(n9581), .D(n9582), .Q(n9563) );
  NOR40 U5086 ( .A(n9619), .B(n9620), .C(n9621), .D(n9622), .Q(n9603) );
  NOR40 U5087 ( .A(n9639), .B(n9640), .C(n9641), .D(n9642), .Q(n9623) );
  NOR40 U5088 ( .A(n9685), .B(n9686), .C(n9687), .D(n9688), .Q(n9669) );
  NOR40 U5089 ( .A(n9665), .B(n9666), .C(n9667), .D(n9668), .Q(n9649) );
  NOR40 U5090 ( .A(n9705), .B(n9706), .C(n9707), .D(n9708), .Q(n9689) );
  NOR40 U5091 ( .A(n9725), .B(n9726), .C(n9727), .D(n9728), .Q(n9709) );
  NOR40 U5092 ( .A(n9769), .B(n9770), .C(n9771), .D(n9772), .Q(n9753) );
  NOR40 U5093 ( .A(n9749), .B(n9750), .C(n9751), .D(n9752), .Q(n9733) );
  NOR40 U5094 ( .A(n9789), .B(n9790), .C(n9791), .D(n9792), .Q(n9773) );
  NOR40 U5095 ( .A(n9809), .B(n9810), .C(n9811), .D(n9812), .Q(n9793) );
  NOR40 U5096 ( .A(n9855), .B(n9856), .C(n9857), .D(n9858), .Q(n9839) );
  NOR40 U5097 ( .A(n9835), .B(n9836), .C(n9837), .D(n9838), .Q(n9819) );
  NOR40 U5098 ( .A(n9875), .B(n9876), .C(n9877), .D(n9878), .Q(n9859) );
  NOR40 U5099 ( .A(n9895), .B(n9896), .C(n9897), .D(n9898), .Q(n9879) );
  NOR40 U5100 ( .A(n9939), .B(n9940), .C(n9941), .D(n9942), .Q(n9923) );
  NOR40 U5101 ( .A(n9919), .B(n9920), .C(n9921), .D(n9922), .Q(n9903) );
  NOR40 U5102 ( .A(n9959), .B(n9960), .C(n9961), .D(n9962), .Q(n9943) );
  NOR40 U5103 ( .A(n9979), .B(n9980), .C(n9981), .D(n9982), .Q(n9963) );
  NOR40 U5104 ( .A(n10025), .B(n10026), .C(n10027), .D(n10028), .Q(n10009) );
  NOR40 U5105 ( .A(n10005), .B(n10006), .C(n10007), .D(n10008), .Q(n9989) );
  NOR40 U5106 ( .A(n10045), .B(n10046), .C(n10047), .D(n10048), .Q(n10029) );
  NOR40 U5107 ( .A(n10065), .B(n10066), .C(n10067), .D(n10068), .Q(n10049) );
  NOR40 U5108 ( .A(n10109), .B(n10110), .C(n10111), .D(n10112), .Q(n10093) );
  NOR40 U5109 ( .A(n10089), .B(n10090), .C(n10091), .D(n10092), .Q(n10073) );
  NOR40 U5110 ( .A(n10129), .B(n10130), .C(n10131), .D(n10132), .Q(n10113) );
  NOR40 U5111 ( .A(n10149), .B(n10150), .C(n10151), .D(n10152), .Q(n10133) );
  NOR40 U5112 ( .A(n10195), .B(n10196), .C(n10197), .D(n10198), .Q(n10179) );
  NOR40 U5113 ( .A(n10175), .B(n10176), .C(n10177), .D(n10178), .Q(n10159) );
  NOR40 U5114 ( .A(n10215), .B(n10216), .C(n10217), .D(n10218), .Q(n10199) );
  NOR40 U5115 ( .A(n10235), .B(n10236), .C(n10237), .D(n10238), .Q(n10219) );
  NOR40 U5116 ( .A(n10279), .B(n10280), .C(n10281), .D(n10282), .Q(n10263) );
  NOR40 U5117 ( .A(n10259), .B(n10260), .C(n10261), .D(n10262), .Q(n10243) );
  NOR40 U5118 ( .A(n10299), .B(n10300), .C(n10301), .D(n10302), .Q(n10283) );
  NOR40 U5119 ( .A(n10319), .B(n10320), .C(n10321), .D(n10322), .Q(n10303) );
  NOR40 U5120 ( .A(n10365), .B(n10366), .C(n10367), .D(n10368), .Q(n10349) );
  NOR40 U5121 ( .A(n10345), .B(n10346), .C(n10347), .D(n10348), .Q(n10329) );
  NOR40 U5122 ( .A(n10385), .B(n10386), .C(n10387), .D(n10388), .Q(n10369) );
  NOR40 U5123 ( .A(n10405), .B(n10406), .C(n10407), .D(n10408), .Q(n10389) );
  NOR40 U5124 ( .A(n10449), .B(n10450), .C(n10451), .D(n10452), .Q(n10433) );
  NOR40 U5125 ( .A(n10429), .B(n10430), .C(n10431), .D(n10432), .Q(n10413) );
  NOR40 U5126 ( .A(n10469), .B(n10470), .C(n10471), .D(n10472), .Q(n10453) );
  NOR40 U5127 ( .A(n10489), .B(n10490), .C(n10491), .D(n10492), .Q(n10473) );
  NOR40 U5128 ( .A(n10535), .B(n10536), .C(n10537), .D(n10538), .Q(n10519) );
  NOR40 U5129 ( .A(n10515), .B(n10516), .C(n10517), .D(n10518), .Q(n10499) );
  NOR40 U5130 ( .A(n10555), .B(n10556), .C(n10557), .D(n10558), .Q(n10539) );
  NOR40 U5131 ( .A(n10575), .B(n10576), .C(n10577), .D(n10578), .Q(n10559) );
  NOR40 U5132 ( .A(n10619), .B(n10620), .C(n10621), .D(n10622), .Q(n10603) );
  NOR40 U5133 ( .A(n10599), .B(n10600), .C(n10601), .D(n10602), .Q(n10583) );
  NOR40 U5134 ( .A(n10639), .B(n10640), .C(n10641), .D(n10642), .Q(n10623) );
  NOR40 U5135 ( .A(n10659), .B(n10660), .C(n10661), .D(n10662), .Q(n10643) );
  NOR40 U5136 ( .A(n10710), .B(n10711), .C(n10712), .D(n10713), .Q(n10692) );
  NOR40 U5137 ( .A(n10688), .B(n10689), .C(n10690), .D(n10691), .Q(n10669) );
  NOR40 U5138 ( .A(n10734), .B(n10735), .C(n10736), .D(n10737), .Q(n10716) );
  NOR40 U5139 ( .A(n10757), .B(n10758), .C(n10759), .D(n10760), .Q(n10740) );
  NOR40 U5140 ( .A(n10806), .B(n10807), .C(n10808), .D(n10809), .Q(n10789) );
  NOR40 U5141 ( .A(n10784), .B(n10785), .C(n10786), .D(n10787), .Q(n10766) );
  NOR40 U5142 ( .A(n10829), .B(n10830), .C(n10831), .D(n10832), .Q(n10811) );
  NOR40 U5143 ( .A(n10867), .B(n10868), .C(n10869), .D(n10870), .Q(n10834) );
  NOR40 U5144 ( .A(n6899), .B(n6900), .C(n6901), .D(n6902), .Q(n6872) );
  NOR40 U5145 ( .A(n7085), .B(n7086), .C(n7087), .D(n7088), .Q(n7074) );
  NOR40 U5146 ( .A(n7255), .B(n7256), .C(n7257), .D(n7258), .Q(n7244) );
  NOR40 U5147 ( .A(n7425), .B(n7426), .C(n7427), .D(n7428), .Q(n7414) );
  NOR40 U5148 ( .A(n7595), .B(n7596), .C(n7597), .D(n7598), .Q(n7584) );
  NOR40 U5149 ( .A(n7765), .B(n7766), .C(n7767), .D(n7768), .Q(n7754) );
  NOR40 U5150 ( .A(n7935), .B(n7936), .C(n7937), .D(n7938), .Q(n7924) );
  NOR40 U5151 ( .A(n8105), .B(n8106), .C(n8107), .D(n8108), .Q(n8094) );
  NOR40 U5152 ( .A(n8275), .B(n8276), .C(n8277), .D(n8278), .Q(n8264) );
  NOR40 U5153 ( .A(n8445), .B(n8446), .C(n8447), .D(n8448), .Q(n8434) );
  NOR40 U5154 ( .A(n8615), .B(n8616), .C(n8617), .D(n8618), .Q(n8604) );
  NOR40 U5155 ( .A(n8785), .B(n8786), .C(n8787), .D(n8788), .Q(n8774) );
  NOR40 U5156 ( .A(n8955), .B(n8956), .C(n8957), .D(n8958), .Q(n8944) );
  NOR40 U5157 ( .A(n9125), .B(n9126), .C(n9127), .D(n9128), .Q(n9114) );
  NOR40 U5158 ( .A(n9295), .B(n9296), .C(n9297), .D(n9298), .Q(n9284) );
  NOR40 U5159 ( .A(n9465), .B(n9466), .C(n9467), .D(n9468), .Q(n9454) );
  NOR40 U5160 ( .A(n9635), .B(n9636), .C(n9637), .D(n9638), .Q(n9624) );
  NOR40 U5161 ( .A(n9805), .B(n9806), .C(n9807), .D(n9808), .Q(n9794) );
  NOR40 U5162 ( .A(n9975), .B(n9976), .C(n9977), .D(n9978), .Q(n9964) );
  NOR40 U5163 ( .A(n10145), .B(n10146), .C(n10147), .D(n10148), .Q(n10134) );
  NOR40 U5164 ( .A(n10315), .B(n10316), .C(n10317), .D(n10318), .Q(n10304) );
  NOR40 U5165 ( .A(n10485), .B(n10486), .C(n10487), .D(n10488), .Q(n10474) );
  NOR40 U5166 ( .A(n10655), .B(n10656), .C(n10657), .D(n10658), .Q(n10644) );
  NOR40 U5167 ( .A(n10847), .B(n10848), .C(n10849), .D(n10850), .Q(n10835) );
  NOR40 U5168 ( .A(n6887), .B(n6888), .C(n6889), .D(n6890), .Q(n6873) );
  NOR40 U5169 ( .A(n7081), .B(n7082), .C(n7083), .D(n7084), .Q(n7075) );
  NOR40 U5170 ( .A(n7251), .B(n7252), .C(n7253), .D(n7254), .Q(n7245) );
  NOR40 U5171 ( .A(n7421), .B(n7422), .C(n7423), .D(n7424), .Q(n7415) );
  NOR40 U5172 ( .A(n7591), .B(n7592), .C(n7593), .D(n7594), .Q(n7585) );
  NOR40 U5173 ( .A(n7761), .B(n7762), .C(n7763), .D(n7764), .Q(n7755) );
  NOR40 U5174 ( .A(n7931), .B(n7932), .C(n7933), .D(n7934), .Q(n7925) );
  NOR40 U5175 ( .A(n8101), .B(n8102), .C(n8103), .D(n8104), .Q(n8095) );
  NOR40 U5176 ( .A(n8271), .B(n8272), .C(n8273), .D(n8274), .Q(n8265) );
  NOR40 U5177 ( .A(n8441), .B(n8442), .C(n8443), .D(n8444), .Q(n8435) );
  NOR40 U5178 ( .A(n8611), .B(n8612), .C(n8613), .D(n8614), .Q(n8605) );
  NOR40 U5179 ( .A(n8781), .B(n8782), .C(n8783), .D(n8784), .Q(n8775) );
  NOR40 U5180 ( .A(n8951), .B(n8952), .C(n8953), .D(n8954), .Q(n8945) );
  NOR40 U5181 ( .A(n9121), .B(n9122), .C(n9123), .D(n9124), .Q(n9115) );
  NOR40 U5182 ( .A(n9291), .B(n9292), .C(n9293), .D(n9294), .Q(n9285) );
  NOR40 U5183 ( .A(n9461), .B(n9462), .C(n9463), .D(n9464), .Q(n9455) );
  NOR40 U5184 ( .A(n9631), .B(n9632), .C(n9633), .D(n9634), .Q(n9625) );
  NOR40 U5185 ( .A(n9801), .B(n9802), .C(n9803), .D(n9804), .Q(n9795) );
  NOR40 U5186 ( .A(n9971), .B(n9972), .C(n9973), .D(n9974), .Q(n9965) );
  NOR40 U5187 ( .A(n10141), .B(n10142), .C(n10143), .D(n10144), .Q(n10135) );
  NOR40 U5188 ( .A(n10311), .B(n10312), .C(n10313), .D(n10314), .Q(n10305) );
  NOR40 U5189 ( .A(n10481), .B(n10482), .C(n10483), .D(n10484), .Q(n10475) );
  NOR40 U5190 ( .A(n10651), .B(n10652), .C(n10653), .D(n10654), .Q(n10645) );
  NOR40 U5191 ( .A(n10843), .B(n10844), .C(n10845), .D(n10846), .Q(n10836) );
  NOR40 U5192 ( .A(n6875), .B(n6876), .C(n6877), .D(n6878), .Q(n6874) );
  NOR40 U5193 ( .A(n7077), .B(n7078), .C(n7079), .D(n7080), .Q(n7076) );
  NOR40 U5194 ( .A(n7247), .B(n7248), .C(n7249), .D(n7250), .Q(n7246) );
  NOR40 U5195 ( .A(n7417), .B(n7418), .C(n7419), .D(n7420), .Q(n7416) );
  NOR40 U5196 ( .A(n7587), .B(n7588), .C(n7589), .D(n7590), .Q(n7586) );
  NOR40 U5197 ( .A(n7757), .B(n7758), .C(n7759), .D(n7760), .Q(n7756) );
  NOR40 U5198 ( .A(n7927), .B(n7928), .C(n7929), .D(n7930), .Q(n7926) );
  NOR40 U5199 ( .A(n8097), .B(n8098), .C(n8099), .D(n8100), .Q(n8096) );
  NOR40 U5200 ( .A(n8267), .B(n8268), .C(n8269), .D(n8270), .Q(n8266) );
  NOR40 U5201 ( .A(n8437), .B(n8438), .C(n8439), .D(n8440), .Q(n8436) );
  NOR40 U5202 ( .A(n8607), .B(n8608), .C(n8609), .D(n8610), .Q(n8606) );
  NOR40 U5203 ( .A(n8777), .B(n8778), .C(n8779), .D(n8780), .Q(n8776) );
  NOR40 U5204 ( .A(n8947), .B(n8948), .C(n8949), .D(n8950), .Q(n8946) );
  NOR40 U5205 ( .A(n9117), .B(n9118), .C(n9119), .D(n9120), .Q(n9116) );
  NOR40 U5206 ( .A(n9287), .B(n9288), .C(n9289), .D(n9290), .Q(n9286) );
  NOR40 U5207 ( .A(n9457), .B(n9458), .C(n9459), .D(n9460), .Q(n9456) );
  NOR40 U5208 ( .A(n9627), .B(n9628), .C(n9629), .D(n9630), .Q(n9626) );
  NOR40 U5209 ( .A(n9797), .B(n9798), .C(n9799), .D(n9800), .Q(n9796) );
  NOR40 U5210 ( .A(n9967), .B(n9968), .C(n9969), .D(n9970), .Q(n9966) );
  NOR40 U5211 ( .A(n10137), .B(n10138), .C(n10139), .D(n10140), .Q(n10136) );
  NOR40 U5212 ( .A(n10307), .B(n10308), .C(n10309), .D(n10310), .Q(n10306) );
  NOR40 U5213 ( .A(n10477), .B(n10478), .C(n10479), .D(n10480), .Q(n10476) );
  NOR40 U5214 ( .A(n10647), .B(n10648), .C(n10649), .D(n10650), .Q(n10646) );
  NOR40 U5215 ( .A(n10838), .B(n10839), .C(n10840), .D(n10841), .Q(n10837) );
  NOR21 U5216 ( .A(n11323), .B(raddr_2), .Q(n10852) );
  NOR21 U5217 ( .A(n11343), .B(raddr_6), .Q(n10686) );
  NOR21 U5218 ( .A(n11322), .B(raddr_3), .Q(n10874) );
  NOR21 U5219 ( .A(n11342), .B(raddr_7), .Q(n10828) );
  INV3 U5220 ( .A(raddr_0), .Q(n11312) );
  INV3 U5221 ( .A(raddr_1), .Q(n11321) );
  INV3 U5222 ( .A(raddr_3), .Q(n11323) );
  INV3 U5223 ( .A(raddr_5), .Q(n11341) );
  INV3 U5224 ( .A(raddr_7), .Q(n11343) );
  INV3 U5225 ( .A(raddr_2), .Q(n11322) );
  INV3 U5226 ( .A(raddr_4), .Q(n11332) );
  INV3 U5227 ( .A(raddr_6), .Q(n11342) );
  BUF2 U5228 ( .A(rclk), .Q(n11298) );
  BUF2 U5229 ( .A(rclk), .Q(n11299) );
  BUF2 U5230 ( .A(rclk), .Q(n11300) );
  BUF2 U5231 ( .A(rclk), .Q(n11301) );
  BUF2 U5232 ( .A(rclk), .Q(n11302) );
  BUF2 U5233 ( .A(rclk), .Q(n11303) );
endmodule


module FIFO_DC_DEPTH256_DWIDTH24_DW01_sub_0 ( .A({A_7, A_6, A_5, A_4, A_3, A_2, 
        A_1, A_0}), .B({B_7, B_6, B_5, B_4, B_3, B_2, B_1, B_0}), CI, .DIFF({
        DIFF_7, DIFF_6, DIFF_5, DIFF_4, DIFF_3, DIFF_2, DIFF_1, DIFF_0}), CO
 );
  input A_7, A_6, A_5, A_4, A_3, A_2, A_1, A_0, B_7, B_6, B_5, B_4, B_3, B_2,
         B_1, B_0, CI;
  output DIFF_7, DIFF_6, DIFF_5, DIFF_4, DIFF_3, DIFF_2, DIFF_1, DIFF_0, CO;
  wire   carry_7, carry_6, carry_5, carry_4, carry_3, carry_2, carry_1, n1, n2,
         n3, n4, n5, n6, n7, n8;

  ADD32 U2_6 ( .A(A_6), .B(n6), .CI(carry_6), .CO(carry_7), .S(DIFF_6) );
  ADD32 U2_5 ( .A(A_5), .B(n5), .CI(carry_5), .CO(carry_6), .S(DIFF_5) );
  ADD32 U2_4 ( .A(A_4), .B(n4), .CI(carry_4), .CO(carry_5), .S(DIFF_4) );
  ADD32 U2_3 ( .A(A_3), .B(n3), .CI(carry_3), .CO(carry_4), .S(DIFF_3) );
  ADD32 U2_2 ( .A(A_2), .B(n2), .CI(carry_2), .CO(carry_3), .S(DIFF_2) );
  ADD32 U2_1 ( .A(A_1), .B(n1), .CI(carry_1), .CO(carry_2), .S(DIFF_1) );
  XOR31 U2_7 ( .A(A_7), .B(n7), .C(carry_7), .Q(DIFF_7) );
  INV3 U1 ( .A(B_1), .Q(n1) );
  INV3 U2 ( .A(A_0), .Q(n8) );
  INV3 U3 ( .A(B_3), .Q(n3) );
  INV3 U4 ( .A(B_5), .Q(n5) );
  INV3 U5 ( .A(B_2), .Q(n2) );
  INV3 U6 ( .A(B_4), .Q(n4) );
  INV3 U7 ( .A(B_6), .Q(n6) );
  INV3 U8 ( .A(B_7), .Q(n7) );
  NAND20 U9 ( .A(B_0), .B(n8), .Q(carry_1) );
endmodule


module FIFO_DC_DEPTH256_DWIDTH24_DW01_inc_0 ( .A({A_7, A_6, A_5, A_4, A_3, A_2, 
        A_1, A_0}), .SUM({SUM_7, SUM_6, SUM_5, SUM_4, SUM_3, SUM_2, SUM_1, 
        SUM_0}) );
  input A_7, A_6, A_5, A_4, A_3, A_2, A_1, A_0;
  output SUM_7, SUM_6, SUM_5, SUM_4, SUM_3, SUM_2, SUM_1, SUM_0;
  wire   carry_7, carry_6, carry_5, carry_4, carry_3, carry_2;

  ADD22 U1_1_6 ( .A(A_6), .B(carry_6), .CO(carry_7), .S(SUM_6) );
  ADD22 U1_1_5 ( .A(A_5), .B(carry_5), .CO(carry_6), .S(SUM_5) );
  ADD22 U1_1_4 ( .A(A_4), .B(carry_4), .CO(carry_5), .S(SUM_4) );
  ADD22 U1_1_3 ( .A(A_3), .B(carry_3), .CO(carry_4), .S(SUM_3) );
  ADD22 U1_1_2 ( .A(A_2), .B(carry_2), .CO(carry_3), .S(SUM_2) );
  ADD21 U1_1_1 ( .A(A_1), .B(A_0), .CO(carry_2), .S(SUM_1) );
  INV3 U1 ( .A(A_0), .Q(SUM_0) );
  XOR20 U2 ( .A(carry_7), .B(A_7), .Q(SUM_7) );
endmodule


module FIFO_DC_DEPTH256_DWIDTH24_DW01_inc_1 ( .A({A_7, A_6, A_5, A_4, A_3, A_2, 
        A_1, A_0}), .SUM({SUM_7, SUM_6, SUM_5, SUM_4, SUM_3, SUM_2, SUM_1, 
        SUM_0}) );
  input A_7, A_6, A_5, A_4, A_3, A_2, A_1, A_0;
  output SUM_7, SUM_6, SUM_5, SUM_4, SUM_3, SUM_2, SUM_1, SUM_0;
  wire   carry_7, carry_6, carry_5, carry_4, carry_3, carry_2;

  ADD22 U1_1_6 ( .A(A_6), .B(carry_6), .CO(carry_7), .S(SUM_6) );
  ADD22 U1_1_5 ( .A(A_5), .B(carry_5), .CO(carry_6), .S(SUM_5) );
  ADD22 U1_1_4 ( .A(A_4), .B(carry_4), .CO(carry_5), .S(SUM_4) );
  ADD22 U1_1_3 ( .A(A_3), .B(carry_3), .CO(carry_4), .S(SUM_3) );
  ADD22 U1_1_2 ( .A(A_2), .B(carry_2), .CO(carry_3), .S(SUM_2) );
  ADD22 U1_1_1 ( .A(A_1), .B(A_0), .CO(carry_2), .S(SUM_1) );
  INV3 U1 ( .A(A_0), .Q(SUM_0) );
  XOR20 U2 ( .A(carry_7), .B(A_7), .Q(SUM_7) );
endmodule


module FIFO_DC_DEPTH256_DWIDTH24 ( rclk, wclk, aclr, .D({D_23, D_22, D_21, 
        D_20, D_19, D_18, D_17, D_16, D_15, D_14, D_13, D_12, D_11, D_10, D_9, 
        D_8, D_7, D_6, D_5, D_4, D_3, D_2, D_1, D_0}), wreq, .Q({Q_23, Q_22, 
        Q_21, Q_20, Q_19, Q_18, Q_17, Q_16, Q_15, Q_14, Q_13, Q_12, Q_11, Q_10, 
        Q_9, Q_8, Q_7, Q_6, Q_5, Q_4, Q_3, Q_2, Q_1, Q_0}), rreq, rd_empty, 
        rd_full, wr_empty, wr_full );
  input rclk, wclk, aclr, D_23, D_22, D_21, D_20, D_19, D_18, D_17, D_16, D_15,
         D_14, D_13, D_12, D_11, D_10, D_9, D_8, D_7, D_6, D_5, D_4, D_3, D_2,
         D_1, D_0, wreq, rreq;
  output Q_23, Q_22, Q_21, Q_20, Q_19, Q_18, Q_17, Q_16, Q_15, Q_14, Q_13,
         Q_12, Q_11, Q_10, Q_9, Q_8, Q_7, Q_6, Q_5, Q_4, Q_3, Q_2, Q_1, Q_0,
         rd_empty, rd_full, wr_empty, wr_full;
  wire   rptr_7, rptr_6, rptr_5, rptr_4, rptr_3, rptr_2, rptr_1, rptr_0, N1,
         N2, N3, N4, N5, N6, N7, N8, wptr_7, wptr_6, wptr_5, wptr_4, wptr_3,
         wptr_2, wptr_1, wptr_0, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N19, N20, N21, N22, N23, N24, N25, N26, rempty, rfull, wempty, wfull,
         n2, n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;
  wire   SYNOPSYS_UNCONNECTED__0;

  DFEC3 rptr_reg_0 ( .D(N1), .E(rreq), .C(rclk), .RN(n5), .Q(rptr_0) );
  DFEC3 rptr_reg_2 ( .D(N3), .E(rreq), .C(rclk), .RN(n5), .Q(rptr_2) );
  DFEC3 rptr_reg_3 ( .D(N4), .E(rreq), .C(rclk), .RN(n5), .Q(rptr_3) );
  DFEC3 rptr_reg_4 ( .D(N5), .E(rreq), .C(rclk), .RN(n5), .Q(rptr_4) );
  DFEC3 rptr_reg_5 ( .D(N6), .E(rreq), .C(rclk), .RN(n4), .Q(rptr_5) );
  DFEC3 rptr_reg_6 ( .D(N7), .E(rreq), .C(rclk), .RN(n4), .Q(rptr_6) );
  DFEC3 rptr_reg_7 ( .D(N8), .E(rreq), .C(rclk), .RN(n4), .Q(rptr_7) );
  DFP3 rempty_reg ( .D(N17), .C(rclk), .SN(n3), .Q(rempty) );
  DFC3 rfull_reg ( .D(N26), .C(rclk), .RN(n3), .Q(rfull) );
  DFC3 rd_full_reg ( .D(rfull), .C(rclk), .RN(n3), .Q(rd_full) );
  DFP3 rd_empty_reg ( .D(rempty), .C(rclk), .SN(n3), .Q(rd_empty) );
  DFP3 wempty_reg ( .D(N17), .C(wclk), .SN(n3), .Q(wempty) );
  DFC3 wfull_reg ( .D(N26), .C(wclk), .RN(n3), .Q(wfull) );
  DFC3 wr_full_reg ( .D(wfull), .C(wclk), .RN(n3), .Q(wr_full) );
  DFP3 wr_empty_reg ( .D(wempty), .C(wclk), .SN(n3), .Q(wr_empty) );
  dual_ported_memory_AWIDTH8_DWIDTH24 mem ( .rclk(rclk), .wclk(wclk), .D({D_23, 
        D_22, D_21, D_20, D_19, D_18, D_17, D_16, D_15, D_14, D_13, D_12, D_11, 
        D_10, D_9, D_8, D_7, D_6, D_5, D_4, D_3, D_2, D_1, D_0}), .waddr({
        wptr_7, wptr_6, wptr_5, wptr_4, wptr_3, wptr_2, wptr_1, wptr_0}), 
        .wreq(wreq), .Q({Q_23, Q_22, Q_21, Q_20, Q_19, Q_18, Q_17, Q_16, Q_15, 
        Q_14, Q_13, Q_12, Q_11, Q_10, Q_9, Q_8, Q_7, Q_6, Q_5, Q_4, Q_3, Q_2, 
        Q_1, Q_0}), .raddr({rptr_7, rptr_6, rptr_5, rptr_4, rptr_3, rptr_2, 
        rptr_1, rptr_0}) );
  FIFO_DC_DEPTH256_DWIDTH24_DW01_sub_0 sub_114 ( .A({wptr_7, wptr_6, wptr_5, 
        wptr_4, wptr_3, wptr_2, wptr_1, wptr_0}), .B({rptr_7, rptr_6, rptr_5, 
        rptr_4, rptr_3, rptr_2, rptr_1, rptr_0}), .CI(n2), .DIFF({N25, N24, 
        N23, N22, N21, N20, N19, SYNOPSYS_UNCONNECTED__0}) );
  FIFO_DC_DEPTH256_DWIDTH24_DW01_inc_0 add_101 ( .A({wptr_7, wptr_6, wptr_5, 
        wptr_4, wptr_3, wptr_2, wptr_1, wptr_0}), .SUM({N16, N15, N14, N13, 
        N12, N11, N10, N9}) );
  FIFO_DC_DEPTH256_DWIDTH24_DW01_inc_1 add_89 ( .A({rptr_7, rptr_6, rptr_5, 
        rptr_4, rptr_3, rptr_2, rptr_1, rptr_0}), .SUM({N8, N7, N6, N5, N4, N3, 
        N2, N1}) );
  DFEC1 wptr_reg_7 ( .D(N16), .E(wreq), .C(wclk), .RN(n3), .Q(wptr_7) );
  DFEC3 wptr_reg_1 ( .D(N10), .E(wreq), .C(wclk), .RN(n4), .Q(wptr_1) );
  DFEC3 wptr_reg_2 ( .D(N11), .E(wreq), .C(wclk), .RN(n4), .Q(wptr_2) );
  DFEC3 wptr_reg_3 ( .D(N12), .E(wreq), .C(wclk), .RN(n4), .Q(wptr_3) );
  DFEC3 wptr_reg_4 ( .D(N13), .E(wreq), .C(wclk), .RN(n4), .Q(wptr_4) );
  DFEC3 wptr_reg_6 ( .D(N15), .E(wreq), .C(wclk), .RN(n4), .Q(wptr_6) );
  DFEC3 wptr_reg_5 ( .D(N14), .E(wreq), .C(wclk), .RN(n4), .Q(wptr_5) );
  DFEC3 wptr_reg_0 ( .D(N9), .E(wreq), .C(wclk), .RN(aclr), .Q(wptr_0), .QN(
        n18) );
  DFEC1 rptr_reg_1 ( .D(N2), .E(rreq), .C(rclk), .RN(n5), .Q(rptr_1), .QN(n1)
         );
  BUF2 U3 ( .A(aclr), .Q(n4) );
  BUF2 U4 ( .A(aclr), .Q(n3) );
  BUF2 U5 ( .A(aclr), .Q(n5) );
  INV3 U6 ( .A(n7), .Q(n19) );
  LOGIC0 U7 ( .Q(n2) );
  XNR20 U8 ( .A(wptr_2), .B(rptr_2), .Q(n11) );
  XNR20 U9 ( .A(wptr_7), .B(rptr_7), .Q(n10) );
  NAND20 U10 ( .A(rptr_0), .B(n18), .Q(n6) );
  AOI220 U11 ( .A(n1), .B(n6), .C(n6), .D(wptr_1), .Q(n7) );
  NOR20 U12 ( .A(n18), .B(rptr_0), .Q(n8) );
  OAI220 U13 ( .A(n8), .B(n1), .C(wptr_1), .D(n8), .Q(n9) );
  NAND40 U14 ( .A(n11), .B(n10), .C(n19), .D(n9), .Q(n17) );
  XNR20 U15 ( .A(wptr_6), .B(rptr_6), .Q(n15) );
  XNR20 U16 ( .A(wptr_5), .B(rptr_5), .Q(n14) );
  XNR20 U17 ( .A(wptr_4), .B(rptr_4), .Q(n13) );
  XNR20 U18 ( .A(wptr_3), .B(rptr_3), .Q(n12) );
  NAND40 U19 ( .A(n15), .B(n14), .C(n13), .D(n12), .Q(n16) );
  NOR20 U20 ( .A(n17), .B(n16), .Q(N17) );
  NAND40 U21 ( .A(N22), .B(N21), .C(N25), .D(N24), .Q(n21) );
  NAND30 U22 ( .A(N19), .B(N23), .C(N20), .Q(n20) );
  NOR20 U23 ( .A(n21), .B(n20), .Q(N26) );
endmodule


module VGA ( CLK_I, RST_I, NRESET, INTA_O, .ADR_I({ADR_I_4, ADR_I_3, ADR_I_2}), 
    .SDAT_I({SDAT_I_31, SDAT_I_30, SDAT_I_29, SDAT_I_28, SDAT_I_27, SDAT_I_26, 
        SDAT_I_25, SDAT_I_24, SDAT_I_23, SDAT_I_22, SDAT_I_21, SDAT_I_20, 
        SDAT_I_19, SDAT_I_18, SDAT_I_17, SDAT_I_16, SDAT_I_15, SDAT_I_14, 
        SDAT_I_13, SDAT_I_12, SDAT_I_11, SDAT_I_10, SDAT_I_9, SDAT_I_8, 
        SDAT_I_7, SDAT_I_6, SDAT_I_5, SDAT_I_4, SDAT_I_3, SDAT_I_2, SDAT_I_1, 
        SDAT_I_0}), .SDAT_O({SDAT_O_31, SDAT_O_30, SDAT_O_29, SDAT_O_28, 
        SDAT_O_27, SDAT_O_26, SDAT_O_25, SDAT_O_24, SDAT_O_23, SDAT_O_22, 
        SDAT_O_21, SDAT_O_20, SDAT_O_19, SDAT_O_18, SDAT_O_17, SDAT_O_16, 
        SDAT_O_15, SDAT_O_14, SDAT_O_13, SDAT_O_12, SDAT_O_11, SDAT_O_10, 
        SDAT_O_9, SDAT_O_8, SDAT_O_7, SDAT_O_6, SDAT_O_5, SDAT_O_4, SDAT_O_3, 
        SDAT_O_2, SDAT_O_1, SDAT_O_0}), .SEL_I({SEL_I_3, SEL_I_2, SEL_I_1, 
        SEL_I_0}), WE_I, STB_I, CYC_I, ACK_O, ERR_O, .ADR_O({ADR_O_31, 
        ADR_O_30, ADR_O_29, ADR_O_28, ADR_O_27, ADR_O_26, ADR_O_25, ADR_O_24, 
        ADR_O_23, ADR_O_22, ADR_O_21, ADR_O_20, ADR_O_19, ADR_O_18, ADR_O_17, 
        ADR_O_16, ADR_O_15, ADR_O_14, ADR_O_13, ADR_O_12, ADR_O_11, ADR_O_10, 
        ADR_O_9, ADR_O_8, ADR_O_7, ADR_O_6, ADR_O_5, ADR_O_4, ADR_O_3, ADR_O_2
        }), .MDAT_I({MDAT_I_31, MDAT_I_30, MDAT_I_29, MDAT_I_28, MDAT_I_27, 
        MDAT_I_26, MDAT_I_25, MDAT_I_24, MDAT_I_23, MDAT_I_22, MDAT_I_21, 
        MDAT_I_20, MDAT_I_19, MDAT_I_18, MDAT_I_17, MDAT_I_16, MDAT_I_15, 
        MDAT_I_14, MDAT_I_13, MDAT_I_12, MDAT_I_11, MDAT_I_10, MDAT_I_9, 
        MDAT_I_8, MDAT_I_7, MDAT_I_6, MDAT_I_5, MDAT_I_4, MDAT_I_3, MDAT_I_2, 
        MDAT_I_1, MDAT_I_0}), .SEL_O({SEL_O_3, SEL_O_2, SEL_O_1, SEL_O_0}), 
        WE_O, STB_O, CYC_O, CAB_O, ACK_I, ERR_I, PCLK, HSYNC, VSYNC, CSYNC, 
        BLANK, .R({R_7, R_6, R_5, R_4, R_3, R_2, R_1, R_0}), .G({G_7, G_6, G_5, 
        G_4, G_3, G_2, G_1, G_0}), .B({B_7, B_6, B_5, B_4, B_3, B_2, B_1, B_0}
        ) );
  input CLK_I, RST_I, NRESET, ADR_I_4, ADR_I_3, ADR_I_2, SDAT_I_31, SDAT_I_30,
         SDAT_I_29, SDAT_I_28, SDAT_I_27, SDAT_I_26, SDAT_I_25, SDAT_I_24,
         SDAT_I_23, SDAT_I_22, SDAT_I_21, SDAT_I_20, SDAT_I_19, SDAT_I_18,
         SDAT_I_17, SDAT_I_16, SDAT_I_15, SDAT_I_14, SDAT_I_13, SDAT_I_12,
         SDAT_I_11, SDAT_I_10, SDAT_I_9, SDAT_I_8, SDAT_I_7, SDAT_I_6,
         SDAT_I_5, SDAT_I_4, SDAT_I_3, SDAT_I_2, SDAT_I_1, SDAT_I_0, SEL_I_3,
         SEL_I_2, SEL_I_1, SEL_I_0, WE_I, STB_I, CYC_I, MDAT_I_31, MDAT_I_30,
         MDAT_I_29, MDAT_I_28, MDAT_I_27, MDAT_I_26, MDAT_I_25, MDAT_I_24,
         MDAT_I_23, MDAT_I_22, MDAT_I_21, MDAT_I_20, MDAT_I_19, MDAT_I_18,
         MDAT_I_17, MDAT_I_16, MDAT_I_15, MDAT_I_14, MDAT_I_13, MDAT_I_12,
         MDAT_I_11, MDAT_I_10, MDAT_I_9, MDAT_I_8, MDAT_I_7, MDAT_I_6,
         MDAT_I_5, MDAT_I_4, MDAT_I_3, MDAT_I_2, MDAT_I_1, MDAT_I_0, ACK_I,
         ERR_I, PCLK;
  output INTA_O, SDAT_O_31, SDAT_O_30, SDAT_O_29, SDAT_O_28, SDAT_O_27,
         SDAT_O_26, SDAT_O_25, SDAT_O_24, SDAT_O_23, SDAT_O_22, SDAT_O_21,
         SDAT_O_20, SDAT_O_19, SDAT_O_18, SDAT_O_17, SDAT_O_16, SDAT_O_15,
         SDAT_O_14, SDAT_O_13, SDAT_O_12, SDAT_O_11, SDAT_O_10, SDAT_O_9,
         SDAT_O_8, SDAT_O_7, SDAT_O_6, SDAT_O_5, SDAT_O_4, SDAT_O_3, SDAT_O_2,
         SDAT_O_1, SDAT_O_0, ACK_O, ERR_O, ADR_O_31, ADR_O_30, ADR_O_29,
         ADR_O_28, ADR_O_27, ADR_O_26, ADR_O_25, ADR_O_24, ADR_O_23, ADR_O_22,
         ADR_O_21, ADR_O_20, ADR_O_19, ADR_O_18, ADR_O_17, ADR_O_16, ADR_O_15,
         ADR_O_14, ADR_O_13, ADR_O_12, ADR_O_11, ADR_O_10, ADR_O_9, ADR_O_8,
         ADR_O_7, ADR_O_6, ADR_O_5, ADR_O_4, ADR_O_3, ADR_O_2, SEL_O_3,
         SEL_O_2, SEL_O_1, SEL_O_0, WE_O, STB_O, CYC_O, CAB_O, HSYNC, VSYNC,
         CSYNC, BLANK, R_7, R_6, R_5, R_4, R_3, R_2, R_1, R_0, G_7, G_6, G_5,
         G_4, G_3, G_2, G_1, G_0, B_7, B_6, B_5, B_4, B_3, B_2, B_1, B_0;
  wire   ctrl_bl, ctrl_csl, ctrl_vsl, ctrl_hsl, ctrl_pc, ctrl_cd_1, ctrl_cd_0,
         ctrl_vbl_1, ctrl_vbl_0, ctrl_cbsw, ctrl_vbsw, ctrl_ven, stat_avmp,
         stat_acmp, bsint, hint, vint, luint, sint, Thsync_7, Thsync_6,
         Thsync_5, Thsync_4, Thsync_3, Thsync_2, Thsync_1, Thsync_0, Thgdel_7,
         Thgdel_6, Thgdel_5, Thgdel_4, Thgdel_3, Thgdel_2, Thgdel_1, Thgdel_0,
         Thgate_15, Thgate_14, Thgate_13, Thgate_12, Thgate_11, Thgate_10,
         Thgate_9, Thgate_8, Thgate_7, Thgate_6, Thgate_5, Thgate_4, Thgate_3,
         Thgate_2, Thgate_1, Thgate_0, Thlen_15, Thlen_14, Thlen_13, Thlen_12,
         Thlen_11, Thlen_10, Thlen_9, Thlen_8, Thlen_7, Thlen_6, Thlen_5,
         Thlen_4, Thlen_3, Thlen_2, Thlen_1, Thlen_0, Tvsync_7, Tvsync_6,
         Tvsync_5, Tvsync_4, Tvsync_3, Tvsync_2, Tvsync_1, Tvsync_0, Tvgdel_7,
         Tvgdel_6, Tvgdel_5, Tvgdel_4, Tvgdel_3, Tvgdel_2, Tvgdel_1, Tvgdel_0,
         Tvgate_15, Tvgate_14, Tvgate_13, Tvgate_12, Tvgate_11, Tvgate_10,
         Tvgate_9, Tvgate_8, Tvgate_7, Tvgate_6, Tvgate_5, Tvgate_4, Tvgate_3,
         Tvgate_2, Tvgate_1, Tvgate_0, Tvlen_15, Tvlen_14, Tvlen_13, Tvlen_12,
         Tvlen_11, Tvlen_10, Tvlen_9, Tvlen_8, Tvlen_7, Tvlen_6, Tvlen_5,
         Tvlen_4, Tvlen_3, Tvlen_2, Tvlen_1, Tvlen_0, VBARa_31, VBARa_30,
         VBARa_29, VBARa_28, VBARa_27, VBARa_26, VBARa_25, VBARa_24, VBARa_23,
         VBARa_22, VBARa_21, VBARa_20, VBARa_19, VBARa_18, VBARa_17, VBARa_16,
         VBARa_15, VBARa_14, VBARa_13, VBARa_12, VBARa_11, VBARa_10, VBARa_9,
         VBARa_8, VBARa_7, VBARa_6, VBARa_5, VBARa_4, VBARa_3, VBARa_2,
         VBARb_31, VBARb_30, VBARb_29, VBARb_28, VBARb_27, VBARb_26, VBARb_25,
         VBARb_24, VBARb_23, VBARb_22, VBARb_21, VBARb_20, VBARb_19, VBARb_18,
         VBARb_17, VBARb_16, VBARb_15, VBARb_14, VBARb_13, VBARb_12, VBARb_11,
         VBARb_10, VBARb_9, VBARb_8, VBARb_7, VBARb_6, VBARb_5, VBARb_4,
         VBARb_3, VBARb_2, CBAR_31, CBAR_30, CBAR_29, CBAR_28, CBAR_27,
         CBAR_26, CBAR_25, CBAR_24, CBAR_23, CBAR_22, CBAR_21, CBAR_20,
         CBAR_19, CBAR_18, CBAR_17, CBAR_16, CBAR_15, CBAR_14, CBAR_13,
         CBAR_12, CBAR_11, line_fifo_wreq, line_fifo_d_23, line_fifo_d_22,
         line_fifo_d_21, line_fifo_d_20, line_fifo_d_19, line_fifo_d_18,
         line_fifo_d_17, line_fifo_d_16, line_fifo_d_15, line_fifo_d_14,
         line_fifo_d_13, line_fifo_d_12, line_fifo_d_11, line_fifo_d_10,
         line_fifo_d_9, line_fifo_d_8, line_fifo_d_7, line_fifo_d_6,
         line_fifo_d_5, line_fifo_d_4, line_fifo_d_3, line_fifo_d_2,
         line_fifo_d_1, line_fifo_d_0, line_fifo_full_wr, cgate, ihsync,
         ivsync, icsync, iblank, line_fifo_empty_rd, luint_pclk, sluint, n2,
         n3, n4;

  DF3 luint_reg ( .D(sluint), .C(CLK_I), .Q(luint) );
  DF3 BLANK_reg ( .D(iblank), .C(PCLK), .Q(BLANK) );
  DF3 CSYNC_reg ( .D(icsync), .C(PCLK), .Q(CSYNC) );
  DF3 VSYNC_reg ( .D(ivsync), .C(PCLK), .Q(VSYNC) );
  DF3 HSYNC_reg ( .D(ihsync), .C(PCLK), .Q(HSYNC) );
  DF3 luint_pclk_reg ( .D(n4), .C(PCLK), .Q(luint_pclk) );
  DF3 sluint_reg ( .D(luint_pclk), .C(CLK_I), .Q(sluint) );
  wb_slave u1 ( .CLK_I(CLK_I), .RST_I(RST_I), .NRESET(NRESET), .ADR_I({ADR_I_4, 
        ADR_I_3, ADR_I_2}), .DAT_I({SDAT_I_31, SDAT_I_30, SDAT_I_29, SDAT_I_28, 
        SDAT_I_27, SDAT_I_26, SDAT_I_25, SDAT_I_24, SDAT_I_23, SDAT_I_22, 
        SDAT_I_21, SDAT_I_20, SDAT_I_19, SDAT_I_18, SDAT_I_17, SDAT_I_16, 
        SDAT_I_15, SDAT_I_14, SDAT_I_13, SDAT_I_12, SDAT_I_11, SDAT_I_10, 
        SDAT_I_9, SDAT_I_8, SDAT_I_7, SDAT_I_6, SDAT_I_5, SDAT_I_4, SDAT_I_3, 
        SDAT_I_2, SDAT_I_1, SDAT_I_0}), .DAT_O({SDAT_O_31, SDAT_O_30, 
        SDAT_O_29, SDAT_O_28, SDAT_O_27, SDAT_O_26, SDAT_O_25, SDAT_O_24, 
        SDAT_O_23, SDAT_O_22, SDAT_O_21, SDAT_O_20, SDAT_O_19, SDAT_O_18, 
        SDAT_O_17, SDAT_O_16, SDAT_O_15, SDAT_O_14, SDAT_O_13, SDAT_O_12, 
        SDAT_O_11, SDAT_O_10, SDAT_O_9, SDAT_O_8, SDAT_O_7, SDAT_O_6, SDAT_O_5, 
        SDAT_O_4, SDAT_O_3, SDAT_O_2, SDAT_O_1, SDAT_O_0}), .SEL_I({SEL_I_3, 
        SEL_I_2, SEL_I_1, SEL_I_0}), .WE_I(WE_I), .STB_I(STB_I), .CYC_I(CYC_I), 
        .ACK_O(ACK_O), .ERR_O(ERR_O), .INTA_O(INTA_O), .BL(ctrl_bl), .CSL(
        ctrl_csl), .VSL(ctrl_vsl), .HSL(ctrl_hsl), .PC(ctrl_pc), .CD({
        ctrl_cd_1, ctrl_cd_0}), .VBL({ctrl_vbl_1, ctrl_vbl_0}), .CBSW(
        ctrl_cbsw), .VBSW(ctrl_vbsw), .Ven(ctrl_ven), .AVMP(stat_avmp), .ACMP(
        stat_acmp), .bsint_in(bsint), .hint_in(hint), .vint_in(vint), 
        .luint_in(luint), .sint_in(sint), .Thsync({Thsync_7, Thsync_6, 
        Thsync_5, Thsync_4, Thsync_3, Thsync_2, Thsync_1, Thsync_0}), .Thgdel(
        {Thgdel_7, Thgdel_6, Thgdel_5, Thgdel_4, Thgdel_3, Thgdel_2, Thgdel_1, 
        Thgdel_0}), .Thgate({Thgate_15, Thgate_14, Thgate_13, Thgate_12, 
        Thgate_11, Thgate_10, Thgate_9, Thgate_8, Thgate_7, Thgate_6, Thgate_5, 
        Thgate_4, Thgate_3, Thgate_2, Thgate_1, Thgate_0}), .Thlen({Thlen_15, 
        Thlen_14, Thlen_13, Thlen_12, Thlen_11, Thlen_10, Thlen_9, Thlen_8, 
        Thlen_7, Thlen_6, Thlen_5, Thlen_4, Thlen_3, Thlen_2, Thlen_1, Thlen_0}), .Tvsync({Tvsync_7, Tvsync_6, Tvsync_5, Tvsync_4, Tvsync_3, Tvsync_2, 
        Tvsync_1, Tvsync_0}), .Tvgdel({Tvgdel_7, Tvgdel_6, Tvgdel_5, Tvgdel_4, 
        Tvgdel_3, Tvgdel_2, Tvgdel_1, Tvgdel_0}), .Tvgate({Tvgate_15, 
        Tvgate_14, Tvgate_13, Tvgate_12, Tvgate_11, Tvgate_10, Tvgate_9, 
        Tvgate_8, Tvgate_7, Tvgate_6, Tvgate_5, Tvgate_4, Tvgate_3, Tvgate_2, 
        Tvgate_1, Tvgate_0}), .Tvlen({Tvlen_15, Tvlen_14, Tvlen_13, Tvlen_12, 
        Tvlen_11, Tvlen_10, Tvlen_9, Tvlen_8, Tvlen_7, Tvlen_6, Tvlen_5, 
        Tvlen_4, Tvlen_3, Tvlen_2, Tvlen_1, Tvlen_0}), .VBARa({VBARa_31, 
        VBARa_30, VBARa_29, VBARa_28, VBARa_27, VBARa_26, VBARa_25, VBARa_24, 
        VBARa_23, VBARa_22, VBARa_21, VBARa_20, VBARa_19, VBARa_18, VBARa_17, 
        VBARa_16, VBARa_15, VBARa_14, VBARa_13, VBARa_12, VBARa_11, VBARa_10, 
        VBARa_9, VBARa_8, VBARa_7, VBARa_6, VBARa_5, VBARa_4, VBARa_3, VBARa_2}), .VBARb({VBARb_31, VBARb_30, VBARb_29, VBARb_28, VBARb_27, VBARb_26, 
        VBARb_25, VBARb_24, VBARb_23, VBARb_22, VBARb_21, VBARb_20, VBARb_19, 
        VBARb_18, VBARb_17, VBARb_16, VBARb_15, VBARb_14, VBARb_13, VBARb_12, 
        VBARb_11, VBARb_10, VBARb_9, VBARb_8, VBARb_7, VBARb_6, VBARb_5, 
        VBARb_4, VBARb_3, VBARb_2}), .CBAR({CBAR_31, CBAR_30, CBAR_29, CBAR_28, 
        CBAR_27, CBAR_26, CBAR_25, CBAR_24, CBAR_23, CBAR_22, CBAR_21, CBAR_20, 
        CBAR_19, CBAR_18, CBAR_17, CBAR_16, CBAR_15, CBAR_14, CBAR_13, CBAR_12, 
        CBAR_11}) );
  wb_master u2 ( .CLK_I(CLK_I), .RST_I(RST_I), .nRESET(NRESET), .CYC_O(CYC_O), 
        .STB_O(STB_O), .CAB_O(CAB_O), .WE_O(WE_O), .ADR_O({ADR_O_31, ADR_O_30, 
        ADR_O_29, ADR_O_28, ADR_O_27, ADR_O_26, ADR_O_25, ADR_O_24, ADR_O_23, 
        ADR_O_22, ADR_O_21, ADR_O_20, ADR_O_19, ADR_O_18, ADR_O_17, ADR_O_16, 
        ADR_O_15, ADR_O_14, ADR_O_13, ADR_O_12, ADR_O_11, ADR_O_10, ADR_O_9, 
        ADR_O_8, ADR_O_7, ADR_O_6, ADR_O_5, ADR_O_4, ADR_O_3, ADR_O_2}), 
        .SEL_O({SEL_O_3, SEL_O_2, SEL_O_1, SEL_O_0}), .ACK_I(ACK_I), .ERR_I(
        ERR_I), .DAT_I({MDAT_I_31, MDAT_I_30, MDAT_I_29, MDAT_I_28, MDAT_I_27, 
        MDAT_I_26, MDAT_I_25, MDAT_I_24, MDAT_I_23, MDAT_I_22, MDAT_I_21, 
        MDAT_I_20, MDAT_I_19, MDAT_I_18, MDAT_I_17, MDAT_I_16, MDAT_I_15, 
        MDAT_I_14, MDAT_I_13, MDAT_I_12, MDAT_I_11, MDAT_I_10, MDAT_I_9, 
        MDAT_I_8, MDAT_I_7, MDAT_I_6, MDAT_I_5, MDAT_I_4, MDAT_I_3, MDAT_I_2, 
        MDAT_I_1, MDAT_I_0}), .SINT(sint), .ctrl_Ven(n3), .ctrl_cd({ctrl_cd_1, 
        ctrl_cd_0}), .ctrl_pc(ctrl_pc), .ctrl_vbl({ctrl_vbl_1, ctrl_vbl_0}), 
        .ctrl_vbsw(ctrl_vbsw), .ctrl_cbsw(ctrl_cbsw), .VBAa({VBARa_31, 
        VBARa_30, VBARa_29, VBARa_28, VBARa_27, VBARa_26, VBARa_25, VBARa_24, 
        VBARa_23, VBARa_22, VBARa_21, VBARa_20, VBARa_19, VBARa_18, VBARa_17, 
        VBARa_16, VBARa_15, VBARa_14, VBARa_13, VBARa_12, VBARa_11, VBARa_10, 
        VBARa_9, VBARa_8, VBARa_7, VBARa_6, VBARa_5, VBARa_4, VBARa_3, VBARa_2}), .VBAb({VBARb_31, VBARb_30, VBARb_29, VBARb_28, VBARb_27, VBARb_26, VBARb_25, 
        VBARb_24, VBARb_23, VBARb_22, VBARb_21, VBARb_20, VBARb_19, VBARb_18, 
        VBARb_17, VBARb_16, VBARb_15, VBARb_14, VBARb_13, VBARb_12, VBARb_11, 
        VBARb_10, VBARb_9, VBARb_8, VBARb_7, VBARb_6, VBARb_5, VBARb_4, 
        VBARb_3, VBARb_2}), .CBA({CBAR_31, CBAR_30, CBAR_29, CBAR_28, CBAR_27, 
        CBAR_26, CBAR_25, CBAR_24, CBAR_23, CBAR_22, CBAR_21, CBAR_20, CBAR_19, 
        CBAR_18, CBAR_17, CBAR_16, CBAR_15, CBAR_14, CBAR_13, CBAR_12, CBAR_11}), .Thgate({Thgate_15, Thgate_14, Thgate_13, Thgate_12, Thgate_11, Thgate_10, 
        Thgate_9, Thgate_8, Thgate_7, Thgate_6, Thgate_5, Thgate_4, Thgate_3, 
        Thgate_2, Thgate_1, Thgate_0}), .Tvgate({Tvgate_15, Tvgate_14, 
        Tvgate_13, Tvgate_12, Tvgate_11, Tvgate_10, Tvgate_9, Tvgate_8, 
        Tvgate_7, Tvgate_6, Tvgate_5, Tvgate_4, Tvgate_3, Tvgate_2, Tvgate_1, 
        Tvgate_0}), .stat_AVMP(stat_avmp), .stat_ACMP(stat_acmp), .bs_req(
        bsint), .line_fifo_wreq(line_fifo_wreq), .line_fifo_d({line_fifo_d_23, 
        line_fifo_d_22, line_fifo_d_21, line_fifo_d_20, line_fifo_d_19, 
        line_fifo_d_18, line_fifo_d_17, line_fifo_d_16, line_fifo_d_15, 
        line_fifo_d_14, line_fifo_d_13, line_fifo_d_12, line_fifo_d_11, 
        line_fifo_d_10, line_fifo_d_9, line_fifo_d_8, line_fifo_d_7, 
        line_fifo_d_6, line_fifo_d_5, line_fifo_d_4, line_fifo_d_3, 
        line_fifo_d_2, line_fifo_d_1, line_fifo_d_0}), .line_fifo_full(
        line_fifo_full_wr) );
  Pgen u3 ( .mclk(CLK_I), .pclk(PCLK), .ctrl_Ven(n3), .ctrl_HSyncL(ctrl_hsl), 
        .Thsync({Thsync_7, Thsync_6, Thsync_5, Thsync_4, Thsync_3, Thsync_2, 
        Thsync_1, Thsync_0}), .Thgdel({Thgdel_7, Thgdel_6, Thgdel_5, Thgdel_4, 
        Thgdel_3, Thgdel_2, Thgdel_1, Thgdel_0}), .Thgate({Thgate_15, 
        Thgate_14, Thgate_13, Thgate_12, Thgate_11, Thgate_10, Thgate_9, 
        Thgate_8, Thgate_7, Thgate_6, Thgate_5, Thgate_4, Thgate_3, Thgate_2, 
        Thgate_1, Thgate_0}), .Thlen({Thlen_15, Thlen_14, Thlen_13, Thlen_12, 
        Thlen_11, Thlen_10, Thlen_9, Thlen_8, Thlen_7, Thlen_6, Thlen_5, 
        Thlen_4, Thlen_3, Thlen_2, Thlen_1, Thlen_0}), .ctrl_VSyncL(ctrl_vsl), 
        .Tvsync({Tvsync_7, Tvsync_6, Tvsync_5, Tvsync_4, Tvsync_3, Tvsync_2, 
        Tvsync_1, Tvsync_0}), .Tvgdel({Tvgdel_7, Tvgdel_6, Tvgdel_5, Tvgdel_4, 
        Tvgdel_3, Tvgdel_2, Tvgdel_1, Tvgdel_0}), .Tvgate({Tvgate_15, 
        Tvgate_14, Tvgate_13, Tvgate_12, Tvgate_11, Tvgate_10, Tvgate_9, 
        Tvgate_8, Tvgate_7, Tvgate_6, Tvgate_5, Tvgate_4, Tvgate_3, Tvgate_2, 
        Tvgate_1, Tvgate_0}), .Tvlen({Tvlen_15, Tvlen_14, Tvlen_13, Tvlen_12, 
        Tvlen_11, Tvlen_10, Tvlen_9, Tvlen_8, Tvlen_7, Tvlen_6, Tvlen_5, 
        Tvlen_4, Tvlen_3, Tvlen_2, Tvlen_1, Tvlen_0}), .ctrl_CSyncL(ctrl_csl), 
        .ctrl_BlankL(ctrl_bl), .eoh(hint), .eov(vint), .Gate(cgate), .Hsync(
        ihsync), .Vsync(ivsync), .Csync(icsync), .Blank(iblank) );
  FIFO_DC_DEPTH256_DWIDTH24 u4 ( .rclk(PCLK), .wclk(CLK_I), .aclr(n3), .D({
        line_fifo_d_23, line_fifo_d_22, line_fifo_d_21, line_fifo_d_20, 
        line_fifo_d_19, line_fifo_d_18, line_fifo_d_17, line_fifo_d_16, 
        line_fifo_d_15, line_fifo_d_14, line_fifo_d_13, line_fifo_d_12, 
        line_fifo_d_11, line_fifo_d_10, line_fifo_d_9, line_fifo_d_8, 
        line_fifo_d_7, line_fifo_d_6, line_fifo_d_5, line_fifo_d_4, 
        line_fifo_d_3, line_fifo_d_2, line_fifo_d_1, line_fifo_d_0}), .wreq(
        line_fifo_wreq), .Q({R_7, R_6, R_5, R_4, R_3, R_2, R_1, R_0, G_7, G_6, 
        G_5, G_4, G_3, G_2, G_1, G_0, B_7, B_6, B_5, B_4, B_3, B_2, B_1, B_0}), 
        .rreq(cgate), .rd_empty(line_fifo_empty_rd), .wr_full(
        line_fifo_full_wr) );
  BUF2 U5 ( .A(ctrl_ven), .Q(n3) );
  INV3 U6 ( .A(n2), .Q(n4) );
  NAND22 U7 ( .A(line_fifo_empty_rd), .B(cgate), .Q(n2) );
endmodule

